--##############################################################################
-- This file was generated automatically from '/src/mips_tb2_template.vhdl'.
-- 
--------------------------------------------------------------------------------
-- Simulation test bench TB2 -- not synthesizable.
--
-- Simulates the CPU core connected to a simulated external static RAM and an
-- internal BRAM block through a stub (i.e. empty).
-- BRAM is initialized with the program object code, and SRAM is initialized 
-- with data secions from program. 
-- The makefile for the source samples include targets to build simulation test 
-- benches using this template, use them as usage examples.
--
-- The memory setup is meant to test the basic 'dummy' cache. 
-- 
-- Console output (at addresses compatible to Plasma's) is logged to text file
-- "hw_sim_console_log.txt".
-- IMPORTANT: The code that echoes UART TX data to the simulation console does
-- line buffering; it will not print anything until it gets a CR (0x0d), and
-- will ifnore LFs (0x0a). Bear this in mind if you see no output when you 
-- expect it.
--
-- WARNING: Will only work on Modelsim; uses custom library SignalSpy.
--##############################################################################

library ieee,modelsim_lib;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mips_pkg.all;


use work.mips_pkg.all;

use modelsim_lib.util.all;
use std.textio.all;
use work.txt_util.all;

entity mips_tb2 is
end;


architecture testbench of mips_tb2 is

-------------------------------------------------------------------------------
-- Simulation parameters

-- Master clock period
constant T : time           := 20 ns;
-- Time the UART is unavailable after writing to the TX register
-- WARNING: slite does not simulate this. The logs may be different when > 0.0!
constant SIMULATED_UART_TX_TIME : time := 0.0 us;

-- Simulation length in clock cycles 
-- 2000 is enough for 'hello' sample, 22000 enough for 10 digits of pi
constant SIMULATION_LENGTH : integer := 22000;

-- Simulated external SRAM size in 32-bit words 
constant SRAM_SIZE : integer := 2048;
-- Ext. SRAM address length (memory is 16 bits wide so it needs an extra address bit)
constant SRAM_ADDR_SIZE : integer := log2(SRAM_SIZE)+1;


-- BRAM table and interface signals --------------------------------------------
constant BRAM_SIZE : integer := 2048;
constant BRAM_ADDR_SIZE : integer := 11;
subtype t_bram_address is std_logic_vector(BRAM_ADDR_SIZE-1 downto 0);
-- (this table holds one byte-slice; the RAM will have 4 of these)
type t_bram is array(0 to BRAM_SIZE-1) of std_logic_vector(7 downto 0);

signal bram_rd_addr :       t_bram_address; 
signal bram_wr_addr :       t_bram_address;
signal bram_rd_data :       t_word;
signal bram_wr_data :       t_word;
signal bram_byte_we :       std_logic_vector(3 downto 0);

-- bram0 is LSB, bram3 is MSB
signal bram3 : t_bram := (
    X"3C",X"27",X"3C",X"24",X"3C",X"24",X"3C",X"27",
    X"AC",X"00",X"14",X"24",X"0C",X"00",X"08",X"23",
    X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",
    X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",
    X"AF",X"AF",X"40",X"23",X"AF",X"00",X"AF",X"00",
    X"AF",X"3C",X"8C",X"00",X"8C",X"00",X"00",X"0C",
    X"23",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
    X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
    X"8F",X"8F",X"8F",X"8F",X"8F",X"00",X"03",X"8F",
    X"00",X"03",X"23",X"34",X"03",X"40",X"40",X"03",
    X"40",X"00",X"00",X"3C",X"24",X"8C",X"00",X"AC",
    X"8C",X"00",X"AC",X"8C",X"00",X"AC",X"8C",X"00",
    X"03",X"AC",X"3C",X"37",X"03",X"00",X"AC",X"AC",
    X"AC",X"AC",X"AC",X"AC",X"AC",X"AC",X"AC",X"AC",
    X"AC",X"AC",X"03",X"34",X"8C",X"8C",X"8C",X"8C",
    X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",
    X"00",X"03",X"34",X"00",X"00",X"00",X"03",X"AC",
    X"00",X"03",X"00",X"30",X"3C",X"AC",X"03",X"00",
    X"03",X"00",X"00",X"24",X"3C",X"24",X"24",X"14",
    X"00",X"00",X"24",X"00",X"00",X"00",X"00",X"24",
    X"30",X"AD",X"00",X"00",X"00",X"14",X"00",X"00",
    X"00",X"14",X"00",X"03",X"00",X"27",X"AF",X"3C",
    X"8E",X"24",X"14",X"00",X"00",X"AF",X"3C",X"3C",
    X"8C",X"8F",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",
    X"AF",X"00",X"10",X"AF",X"3C",X"26",X"00",X"00",
    X"00",X"02",X"AE",X"26",X"16",X"00",X"00",X"00",
    X"24",X"00",X"AC",X"3C",X"00",X"3C",X"AE",X"10",
    X"AE",X"3C",X"3C",X"26",X"8E",X"02",X"24",X"24",
    X"00",X"01",X"8D",X"24",X"00",X"24",X"24",X"AE",
    X"AC",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
    X"AD",X"00",X"11",X"AE",X"00",X"02",X"24",X"24",
    X"01",X"8D",X"01",X"25",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"14",X"00",X"00",X"24",X"00",
    X"AD",X"00",X"15",X"25",X"02",X"25",X"00",X"01",
    X"AE",X"AC",X"AE",X"14",X"00",X"00",X"24",X"AF",
    X"AF",X"00",X"0C",X"00",X"8E",X"8E",X"8F",X"14",
    X"00",X"00",X"AE",X"00",X"AE",X"8F",X"00",X"14",
    X"AE",X"8F",X"00",X"8F",X"8F",X"8F",X"8F",X"8F",
    X"8F",X"8F",X"8F",X"8F",X"03",X"27",X"44",X"3C",
    X"00",X"44",X"03",X"00",X"44",X"44",X"00",X"00",
    X"3C",X"34",X"30",X"30",X"00",X"3C",X"00",X"00",
    X"00",X"11",X"00",X"00",X"28",X"11",X"00",X"00",
    X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
    X"00",X"10",X"3C",X"00",X"10",X"3C",X"3C",X"00",
    X"00",X"14",X"24",X"3C",X"00",X"14",X"00",X"3C",
    X"00",X"00",X"10",X"24",X"18",X"3C",X"34",X"00",
    X"00",X"00",X"00",X"00",X"00",X"44",X"03",X"00",
    X"00",X"28",X"11",X"00",X"00",X"08",X"00",X"00",
    X"08",X"00",X"08",X"00",X"00",X"14",X"3C",X"44",
    X"03",X"00",X"00",X"44",X"03",X"00",X"44",X"3C",
    X"00",X"44",X"08",X"00",X"44",X"44",X"3C",X"34",
    X"3C",X"00",X"00",X"00",X"01",X"30",X"31",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
    X"31",X"01",X"00",X"00",X"30",X"00",X"01",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
    X"00",X"10",X"00",X"30",X"00",X"3C",X"24",X"30",
    X"00",X"10",X"00",X"3C",X"00",X"00",X"14",X"24",
    X"18",X"00",X"3C",X"34",X"00",X"00",X"00",X"00",
    X"00",X"00",X"44",X"03",X"00",X"44",X"03",X"00",
    X"00",X"44",X"03",X"00",X"44",X"44",X"3C",X"35",
    X"3C",X"00",X"00",X"00",X"01",X"00",X"00",X"14",
    X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"01",
    X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"31",
    X"01",X"00",X"00",X"31",X"00",X"01",X"01",X"00",
    X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",
    X"01",X"00",X"14",X"00",X"00",X"00",X"00",X"10",
    X"00",X"30",X"00",X"3C",X"24",X"30",X"00",X"10",
    X"00",X"3C",X"00",X"00",X"14",X"24",X"04",X"00",
    X"10",X"00",X"3C",X"34",X"00",X"00",X"00",X"00",
    X"00",X"00",X"44",X"03",X"00",X"44",X"03",X"00",
    X"00",X"44",X"03",X"00",X"44",X"3C",X"34",X"3C",
    X"00",X"00",X"00",X"30",X"24",X"00",X"18",X"00",
    X"28",X"10",X"00",X"00",X"04",X"00",X"00",X"03",
    X"00",X"08",X"00",X"04",X"00",X"10",X"3C",X"00",
    X"10",X"00",X"24",X"3C",X"00",X"00",X"14",X"24",
    X"3C",X"00",X"14",X"3C",X"3C",X"00",X"00",X"10",
    X"24",X"3C",X"34",X"00",X"00",X"00",X"00",X"00",
    X"00",X"44",X"03",X"00",X"00",X"14",X"3C",X"00",
    X"44",X"03",X"00",X"08",X"24",X"44",X"44",X"00",
    X"10",X"00",X"00",X"00",X"00",X"14",X"00",X"14",
    X"00",X"14",X"24",X"24",X"00",X"00",X"30",X"30",
    X"00",X"14",X"00",X"14",X"3C",X"34",X"00",X"00",
    X"3C",X"00",X"00",X"00",X"14",X"00",X"00",X"03",
    X"00",X"03",X"24",X"03",X"24",X"03",X"00",X"08",
    X"00",X"08",X"00",X"08",X"00",X"08",X"00",X"44",
    X"44",X"00",X"00",X"03",X"00",X"44",X"44",X"00",
    X"00",X"03",X"00",X"27",X"24",X"AF",X"AF",X"AF",
    X"AF",X"AF",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",
    X"E7",X"46",X"0C",X"E7",X"46",X"46",X"0C",X"46",
    X"46",X"0C",X"46",X"44",X"0C",X"24",X"46",X"46",
    X"0C",X"46",X"46",X"0C",X"46",X"44",X"00",X"08",
    X"24",X"44",X"46",X"46",X"12",X"26",X"0C",X"46",
    X"44",X"0C",X"46",X"44",X"44",X"0C",X"46",X"46",
    X"0C",X"46",X"46",X"0C",X"46",X"46",X"46",X"0C",
    X"46",X"46",X"0C",X"46",X"02",X"16",X"46",X"46",
    X"C7",X"C7",X"C7",X"C7",X"8F",X"8F",X"8F",X"8F",
    X"8F",X"C7",X"C7",X"C7",X"C7",X"03",X"27",X"27",
    X"3C",X"E7",X"E7",X"E7",X"E7",X"AF",X"AF",X"AF",
    X"AF",X"AF",X"E7",X"E7",X"C4",X"08",X"46",X"0C",
    X"00",X"46",X"46",X"0C",X"46",X"46",X"1C",X"46",
    X"44",X"0C",X"46",X"46",X"04",X"46",X"0C",X"00",
    X"46",X"44",X"0C",X"46",X"46",X"04",X"46",X"3C",
    X"C6",X"0C",X"46",X"04",X"46",X"0C",X"46",X"24",
    X"0C",X"46",X"44",X"3C",X"3C",X"C4",X"0C",X"46",
    X"04",X"00",X"C6",X"0C",X"46",X"3C",X"46",X"00",
    X"46",X"0C",X"46",X"44",X"C6",X"3C",X"02",X"46",
    X"46",X"24",X"24",X"44",X"0C",X"46",X"26",X"00",
    X"46",X"00",X"0C",X"26",X"46",X"0C",X"46",X"46",
    X"46",X"0C",X"46",X"46",X"0C",X"46",X"16",X"46",
    X"C7",X"C7",X"C7",X"44",X"8F",X"8F",X"8F",X"8F",
    X"8F",X"C7",X"C7",X"C7",X"46",X"08",X"27",X"3C",
    X"8E",X"08",X"3C",X"3C",X"C4",X"27",X"AF",X"0C",
    X"00",X"46",X"8F",X"08",X"27",X"44",X"27",X"AF",
    X"AF",X"AF",X"AF",X"E7",X"E7",X"E7",X"44",X"0C",
    X"E7",X"04",X"3C",X"C4",X"44",X"0C",X"46",X"1C",
    X"3C",X"C4",X"44",X"0C",X"00",X"18",X"3C",X"C4",
    X"44",X"0C",X"46",X"44",X"46",X"0C",X"46",X"3C",
    X"C4",X"0C",X"46",X"46",X"0C",X"46",X"0C",X"46",
    X"3C",X"C4",X"0C",X"46",X"3C",X"C4",X"46",X"C7",
    X"C7",X"8F",X"8F",X"8F",X"8F",X"C7",X"C7",X"08",
    X"27",X"44",X"0C",X"46",X"0C",X"46",X"3C",X"C4",
    X"08",X"46",X"3C",X"C4",X"44",X"0C",X"00",X"04",
    X"3C",X"02",X"44",X"44",X"44",X"0C",X"02",X"46",
    X"24",X"24",X"46",X"0C",X"46",X"02",X"0C",X"46",
    X"46",X"0C",X"46",X"44",X"0C",X"46",X"26",X"44",
    X"16",X"46",X"C7",X"C7",X"8F",X"44",X"8F",X"8F",
    X"8F",X"C7",X"C7",X"03",X"27",X"3C",X"C4",X"44",
    X"0C",X"00",X"18",X"3C",X"3C",X"C4",X"44",X"0C",
    X"00",X"0C",X"46",X"3C",X"C4",X"08",X"46",X"3C",
    X"3C",X"C4",X"02",X"44",X"0C",X"46",X"44",X"46",
    X"0C",X"46",X"3C",X"C4",X"0C",X"46",X"46",X"0C",
    X"46",X"0C",X"46",X"3C",X"C4",X"0C",X"46",X"3C",
    X"C4",X"0C",X"46",X"44",X"08",X"02",X"27",X"AF",
    X"E7",X"E7",X"E7",X"46",X"E7",X"0C",X"46",X"0C",
    X"46",X"44",X"46",X"0C",X"E7",X"C7",X"04",X"00",
    X"C7",X"C7",X"8F",X"C7",X"C7",X"03",X"27",X"44",
    X"0C",X"46",X"C7",X"18",X"3C",X"C7",X"C7",X"C4",
    X"8F",X"C7",X"C7",X"46",X"08",X"27",X"C7",X"C7",
    X"C4",X"8F",X"C7",X"C7",X"46",X"08",X"27",X"27",
    X"3C",X"AF",X"AF",X"E7",X"E7",X"3C",X"3C",X"C4",
    X"3C",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",X"E7",
    X"E7",X"AF",X"C4",X"C6",X"C6",X"08",X"46",X"0C",
    X"00",X"46",X"46",X"0C",X"46",X"46",X"46",X"0C",
    X"46",X"46",X"1C",X"46",X"3C",X"C6",X"C4",X"08",
    X"46",X"0C",X"00",X"46",X"46",X"0C",X"46",X"46",
    X"46",X"0C",X"46",X"46",X"04",X"46",X"C6",X"46",
    X"0C",X"46",X"46",X"46",X"24",X"24",X"46",X"0C",
    X"46",X"02",X"0C",X"46",X"46",X"0C",X"46",X"46",
    X"46",X"0C",X"46",X"46",X"0C",X"46",X"26",X"16",
    X"46",X"C7",X"C7",X"C7",X"C7",X"46",X"C7",X"8F",
    X"8F",X"8F",X"C7",X"C7",X"C7",X"C7",X"C7",X"46",
    X"08",X"27",X"27",X"3C",X"E7",X"E7",X"C4",X"3C",
    X"E7",X"E7",X"C4",X"3C",X"E7",X"E7",X"E7",X"E7",
    X"E7",X"E7",X"AF",X"AF",X"AF",X"AF",X"C4",X"44",
    X"08",X"46",X"0C",X"00",X"46",X"46",X"0C",X"46",
    X"46",X"46",X"0C",X"46",X"46",X"1C",X"46",X"3C",
    X"3C",X"C4",X"3C",X"C4",X"C6",X"08",X"00",X"0C",
    X"00",X"46",X"46",X"0C",X"46",X"46",X"46",X"0C",
    X"46",X"46",X"1C",X"46",X"3C",X"C4",X"3C",X"C6",
    X"C4",X"08",X"00",X"0C",X"00",X"46",X"46",X"0C",
    X"46",X"46",X"46",X"0C",X"46",X"46",X"04",X"46",
    X"3C",X"C4",X"0C",X"3C",X"44",X"3C",X"C4",X"44",
    X"02",X"24",X"24",X"44",X"0C",X"46",X"02",X"0C",
    X"46",X"46",X"0C",X"46",X"46",X"0C",X"46",X"26",
    X"16",X"46",X"C7",X"C7",X"C7",X"C7",X"46",X"C7",
    X"8F",X"8F",X"8F",X"8F",X"C7",X"C7",X"C7",X"C7",
    X"C7",X"46",X"08",X"27",X"27",X"AF",X"0C",X"E7",
    X"C7",X"00",X"46",X"0C",X"46",X"46",X"8F",X"08",
    X"27",X"10",X"00",X"30",X"10",X"00",X"00",X"14",
    X"00",X"03",X"00",X"00",X"00",X"00",X"08",X"24",
    X"10",X"01",X"00",X"30",X"00",X"24",X"00",X"00",
    X"15",X"00",X"10",X"2C",X"11",X"00",X"00",X"34",
    X"14",X"01",X"03",X"00",X"04",X"00",X"04",X"00",
    X"00",X"00",X"00",X"08",X"24",X"10",X"01",X"00",
    X"30",X"00",X"24",X"00",X"00",X"15",X"00",X"10",
    X"2C",X"11",X"00",X"00",X"34",X"14",X"01",X"11",
    X"00",X"00",X"03",X"00",X"00",X"04",X"24",X"00",
    X"08",X"39",X"00",X"00",X"00",X"08",X"24",X"10",
    X"01",X"00",X"30",X"00",X"24",X"00",X"15",X"00",
    X"10",X"2C",X"11",X"00",X"00",X"14",X"01",X"03",
    X"00",X"00",X"00",X"00",X"08",X"24",X"10",X"01",
    X"00",X"30",X"00",X"24",X"00",X"15",X"00",X"10",
    X"2C",X"11",X"00",X"00",X"14",X"01",X"03",X"00",
    X"40",X"40",X"3F",X"3F",X"BF",X"BF",X"3E",X"3E",
    X"3E",X"3D",X"BE",X"40",X"C0",X"40",X"3E",X"3D",
    X"40",X"41",X"3F",X"3F",X"3F",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal bram2 : t_bram := (
    X"1C",X"9C",X"05",X"A5",X"04",X"84",X"1D",X"BD",
    X"A0",X"A4",X"60",X"A5",X"00",X"00",X"00",X"BD",
    X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",
    X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B8",
    X"B9",X"BF",X"1A",X"5A",X"BA",X"00",X"BB",X"00",
    X"BB",X"06",X"C4",X"00",X"C6",X"00",X"86",X"00",
    X"A5",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",
    X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",
    X"B8",X"B9",X"BF",X"BA",X"BB",X"00",X"60",X"BB",
    X"00",X"60",X"BD",X"1B",X"40",X"9B",X"02",X"E0",
    X"84",X"00",X"00",X"05",X"A5",X"A6",X"00",X"06",
    X"A6",X"00",X"06",X"A6",X"00",X"06",X"A6",X"00",
    X"E0",X"06",X"1A",X"5A",X"40",X"00",X"90",X"91",
    X"92",X"93",X"94",X"95",X"96",X"97",X"9E",X"9C",
    X"9D",X"9F",X"E0",X"02",X"90",X"91",X"92",X"93",
    X"94",X"95",X"96",X"97",X"9E",X"9C",X"9D",X"9F",
    X"00",X"E0",X"A2",X"85",X"00",X"00",X"E0",X"C4",
    X"00",X"E0",X"00",X"84",X"02",X"44",X"E0",X"00",
    X"E0",X"00",X"00",X"02",X"08",X"06",X"07",X"40",
    X"82",X"07",X"63",X"00",X"00",X"00",X"A2",X"A5",
    X"A5",X"05",X"00",X"00",X"00",X"C0",X"46",X"07",
    X"00",X"67",X"85",X"E0",X"00",X"BD",X"B2",X"12",
    X"43",X"06",X"C0",X"66",X"07",X"BE",X"02",X"1E",
    X"47",X"C5",X"BF",X"B7",X"B6",X"B5",X"B4",X"B3",
    X"B1",X"00",X"E5",X"B0",X"10",X"10",X"07",X"05",
    X"90",X"08",X"06",X"10",X"04",X"00",X"07",X"A4",
    X"E7",X"E4",X"47",X"16",X"05",X"17",X"C0",X"C0",
    X"E6",X"11",X"10",X"10",X"27",X"00",X"15",X"13",
    X"05",X"10",X"04",X"C9",X"64",X"CC",X"AA",X"EC",
    X"4A",X"00",X"00",X"00",X"20",X"89",X"07",X"00",
    X"09",X"00",X"40",X"C4",X"0A",X"89",X"C6",X"A8",
    X"44",X"2B",X"00",X"08",X"00",X"00",X"00",X"6B",
    X"00",X"8B",X"00",X"C0",X"86",X"07",X"C6",X"00",
    X"2B",X"00",X"15",X"29",X"65",X"8C",X"06",X"86",
    X"EC",X"40",X"C4",X"60",X"83",X"07",X"A5",X"C5",
    X"A2",X"00",X"00",X"87",X"C7",X"43",X"C5",X"60",
    X"E3",X"07",X"C0",X"05",X"E6",X"A2",X"00",X"C0",
    X"27",X"BF",X"00",X"BE",X"B7",X"B6",X"B5",X"B4",
    X"B3",X"B2",X"B1",X"B0",X"E0",X"BD",X"02",X"03",
    X"62",X"82",X"E0",X"00",X"04",X"02",X"04",X"02",
    X"05",X"A5",X"63",X"E7",X"45",X"08",X"85",X"E3",
    X"C8",X"20",X"A8",X"67",X"E8",X"00",X"00",X"E6",
    X"81",X"00",X"05",X"41",X"00",X"06",X"C5",X"C0",
    X"C0",X"40",X"04",X"44",X"80",X"04",X"05",X"02",
    X"45",X"80",X"63",X"04",X"44",X"80",X"00",X"05",
    X"02",X"45",X"80",X"63",X"60",X"04",X"84",X"06",
    X"44",X"06",X"46",X"03",X"43",X"83",X"E0",X"00",
    X"E3",X"68",X"00",X"00",X"65",X"00",X"E0",X"E0",
    X"00",X"00",X"00",X"00",X"06",X"40",X"04",X"80",
    X"E0",X"00",X"00",X"83",X"E0",X"00",X"03",X"02",
    X"62",X"82",X"00",X"00",X"07",X"06",X"05",X"A5",
    X"02",X"C5",X"E5",X"A2",X"02",X"A4",X"02",X"44",
    X"05",X"08",X"00",X"09",X"00",X"45",X"00",X"22",
    X"23",X"04",X"09",X"00",X"82",X"04",X"05",X"62",
    X"03",X"03",X"02",X"00",X"85",X"89",X"2A",X"09",
    X"49",X"40",X"07",X"A5",X"06",X"04",X"A5",X"63",
    X"44",X"80",X"A3",X"05",X"02",X"45",X"80",X"63",
    X"60",X"E6",X"04",X"84",X"06",X"44",X"06",X"46",
    X"03",X"43",X"83",X"E0",X"00",X"80",X"E0",X"00",
    X"00",X"83",X"E0",X"00",X"07",X"06",X"08",X"08",
    X"03",X"C8",X"E8",X"A3",X"03",X"08",X"05",X"60",
    X"83",X"07",X"AB",X"05",X"00",X"04",X"89",X"2B",
    X"04",X"00",X"02",X"00",X"4B",X"00",X"4B",X"6C",
    X"25",X"0B",X"00",X"22",X"09",X"45",X"82",X"02",
    X"02",X"02",X"00",X"25",X"AB",X"6C",X"0B",X"4B",
    X"02",X"02",X"60",X"43",X"07",X"00",X"44",X"40",
    X"07",X"A5",X"06",X"04",X"A5",X"63",X"44",X"80",
    X"A3",X"05",X"02",X"45",X"80",X"63",X"60",X"00",
    X"60",X"E6",X"04",X"84",X"06",X"44",X"06",X"46",
    X"03",X"43",X"83",X"E0",X"00",X"80",X"E0",X"00",
    X"00",X"83",X"E0",X"00",X"03",X"02",X"42",X"05",
    X"03",X"62",X"45",X"84",X"05",X"A4",X"80",X"02",
    X"85",X"A0",X"00",X"82",X"61",X"00",X"02",X"E0",
    X"00",X"00",X"00",X"80",X"80",X"40",X"03",X"43",
    X"60",X"00",X"03",X"06",X"02",X"46",X"A0",X"63",
    X"05",X"45",X"A0",X"05",X"06",X"02",X"46",X"A0",
    X"63",X"05",X"A5",X"45",X"03",X"04",X"62",X"04",
    X"44",X"82",X"E0",X"00",X"04",X"40",X"03",X"00",
    X"82",X"E0",X"00",X"00",X"03",X"03",X"04",X"00",
    X"64",X"00",X"03",X"04",X"A2",X"C0",X"45",X"A0",
    X"00",X"40",X"02",X"02",X"03",X"04",X"C6",X"A5",
    X"A6",X"E0",X"C5",X"A0",X"05",X"A5",X"85",X"65",
    X"05",X"85",X"65",X"85",X"A0",X"00",X"02",X"E0",
    X"00",X"E0",X"02",X"E0",X"02",X"E0",X"02",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
    X"02",X"00",X"62",X"E0",X"02",X"03",X"02",X"00",
    X"62",X"E0",X"02",X"BD",X"04",X"BF",X"B3",X"B2",
    X"B1",X"B0",X"BA",X"BB",X"B6",X"B7",X"B4",X"B5",
    X"B8",X"00",X"00",X"B9",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"11",X"00",X"04",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
    X"12",X"10",X"00",X"00",X"30",X"73",X"00",X"00",
    X"90",X"00",X"00",X"91",X"90",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"72",X"00",X"00",
    X"BA",X"B8",X"B6",X"B4",X"BF",X"B3",X"B2",X"B1",
    X"B0",X"BB",X"B9",X"B7",X"B5",X"E0",X"BD",X"BD",
    X"02",X"B6",X"B7",X"B4",X"B5",X"BF",X"B3",X"B2",
    X"B1",X"B0",X"B8",X"B9",X"54",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
    X"80",X"00",X"00",X"00",X"41",X"00",X"00",X"00",
    X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"10",
    X"14",X"00",X"00",X"40",X"00",X"00",X"00",X"04",
    X"00",X"00",X"11",X"12",X"02",X"4E",X"00",X"00",
    X"40",X"00",X"0C",X"00",X"00",X"02",X"00",X"51",
    X"00",X"00",X"00",X"02",X"54",X"13",X"62",X"00",
    X"00",X"12",X"10",X"93",X"00",X"00",X"44",X"92",
    X"00",X"00",X"00",X"52",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
    X"B8",X"B6",X"B4",X"91",X"BF",X"B3",X"B2",X"B1",
    X"B0",X"B9",X"B7",X"B5",X"00",X"00",X"BD",X"12",
    X"51",X"00",X"02",X"02",X"4E",X"BD",X"BF",X"00",
    X"00",X"00",X"BF",X"00",X"BD",X"80",X"BD",X"B0",
    X"BF",X"B2",X"B1",X"B6",X"B7",X"B4",X"10",X"00",
    X"B5",X"40",X"02",X"54",X"90",X"00",X"00",X"40",
    X"02",X"4E",X"90",X"00",X"00",X"40",X"02",X"54",
    X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"02",
    X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"02",X"4C",X"00",X"00",X"02",X"4E",X"00",X"B6",
    X"B4",X"BF",X"B2",X"B1",X"B0",X"B7",X"B5",X"00",
    X"BD",X"90",X"00",X"00",X"00",X"00",X"02",X"4C",
    X"00",X"00",X"02",X"4E",X"90",X"00",X"00",X"40",
    X"02",X"02",X"90",X"82",X"90",X"00",X"00",X"00",
    X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"92",X"00",X"00",X"10",X"12",
    X"11",X"00",X"B6",X"B4",X"BF",X"92",X"B2",X"B1",
    X"B0",X"B7",X"B5",X"E0",X"BD",X"02",X"4E",X"90",
    X"00",X"00",X"40",X"02",X"02",X"4C",X"90",X"00",
    X"00",X"00",X"00",X"02",X"4C",X"00",X"00",X"02",
    X"11",X"54",X"30",X"90",X"00",X"00",X"90",X"00",
    X"00",X"00",X"02",X"4C",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"02",X"4C",X"00",X"00",X"02",
    X"4E",X"00",X"00",X"12",X"00",X"32",X"BD",X"BF",
    X"B6",X"B7",X"B4",X"00",X"B5",X"00",X"00",X"00",
    X"00",X"80",X"00",X"00",X"A0",X"A0",X"40",X"00",
    X"B6",X"B4",X"BF",X"B7",X"B5",X"E0",X"BD",X"80",
    X"00",X"00",X"A0",X"40",X"02",X"B6",X"B4",X"4E",
    X"BF",X"B7",X"B5",X"00",X"00",X"BD",X"B6",X"B4",
    X"4E",X"BF",X"B7",X"B5",X"00",X"00",X"BD",X"BD",
    X"02",X"B1",X"B0",X"B8",X"B9",X"10",X"11",X"58",
    X"02",X"BC",X"BD",X"BA",X"BB",X"B6",X"B7",X"B4",
    X"B5",X"BF",X"5A",X"16",X"3C",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"40",X"00",X"02",X"3A",X"5C",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"40",X"00",X"18",X"00",
    X"00",X"00",X"00",X"00",X"10",X"11",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",
    X"00",X"BC",X"BA",X"B8",X"B4",X"00",X"B6",X"BF",
    X"B1",X"B0",X"BD",X"BB",X"B9",X"B7",X"B5",X"00",
    X"00",X"BD",X"BD",X"02",X"B8",X"B9",X"58",X"02",
    X"BA",X"BB",X"5A",X"02",X"BC",X"BD",X"B6",X"B7",
    X"B4",X"B5",X"BF",X"B2",X"B1",X"B0",X"5C",X"80",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"02",
    X"10",X"58",X"02",X"5C",X"1A",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"40",X"00",X"02",X"5A",X"02",X"18",
    X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
    X"02",X"4E",X"00",X"12",X"02",X"03",X"74",X"80",
    X"42",X"10",X"11",X"92",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
    X"11",X"00",X"BC",X"BA",X"B8",X"B4",X"00",X"B6",
    X"BF",X"B2",X"B1",X"B0",X"BD",X"BB",X"B9",X"B7",
    X"B5",X"00",X"00",X"BD",X"BD",X"BF",X"00",X"AE",
    X"AE",X"00",X"00",X"00",X"00",X"00",X"BF",X"00",
    X"BD",X"A0",X"00",X"A3",X"60",X"05",X"44",X"A0",
    X"04",X"E0",X"00",X"05",X"00",X"00",X"00",X"0A",
    X"CA",X"07",X"05",X"A8",X"83",X"C6",X"03",X"08",
    X"20",X"02",X"60",X"A9",X"20",X"00",X"83",X"42",
    X"CA",X"07",X"E0",X"00",X"80",X"00",X"A0",X"00",
    X"05",X"00",X"00",X"00",X"0A",X"CA",X"07",X"05",
    X"A8",X"83",X"C6",X"03",X"08",X"20",X"02",X"60",
    X"A9",X"20",X"00",X"83",X"42",X"CA",X"07",X"60",
    X"00",X"02",X"E0",X"00",X"04",X"A1",X"0B",X"05",
    X"00",X"6B",X"80",X"05",X"00",X"00",X"04",X"C4",
    X"07",X"05",X"A8",X"43",X"C6",X"03",X"20",X"08",
    X"60",X"A9",X"20",X"00",X"43",X"C4",X"07",X"E0",
    X"00",X"80",X"05",X"00",X"00",X"04",X"C4",X"07",
    X"05",X"A8",X"43",X"C6",X"03",X"20",X"08",X"60",
    X"A9",X"20",X"00",X"43",X"C4",X"07",X"E0",X"00",
    X"C9",X"49",X"80",X"C9",X"80",X"C9",X"E6",X"BF",
    X"C9",X"0D",X"E6",X"EC",X"00",X"00",X"0A",X"80",
    X"31",X"80",X"00",X"31",X"C0",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal bram1 : t_bram := (
    X"80",X"80",X"80",X"00",X"80",X"03",X"80",X"02",
    X"00",X"18",X"FF",X"00",X"00",X"00",X"00",X"FF",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"70",X"FF",X"00",X"D8",X"00",X"D8",
    X"00",X"20",X"00",X"00",X"00",X"00",X"20",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"00",
    X"60",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"10",X"20",X"00",X"00",
    X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"10",
    X"00",X"00",X"18",X"03",X"20",X"00",X"00",X"00",
    X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"00",
    X"00",X"00",X"28",X"00",X"00",X"00",X"00",X"00",
    X"10",X"FF",X"20",X"00",X"00",X"FF",X"00",X"80",
    X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"30",X"00",X"00",X"80",X"02",X"40",X"20",
    X"20",X"80",X"00",X"00",X"FF",X"00",X"20",X"20",
    X"00",X"38",X"00",X"80",X"30",X"80",X"00",X"00",
    X"00",X"80",X"80",X"02",X"00",X"A0",X"FF",X"00",
    X"40",X"40",X"00",X"FF",X"00",X"FF",X"FF",X"00",
    X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"48",
    X"00",X"20",X"00",X"00",X"48",X"48",X"FF",X"FF",
    X"00",X"00",X"50",X"FF",X"20",X"00",X"00",X"00",
    X"58",X"20",X"00",X"00",X"00",X"00",X"FF",X"58",
    X"00",X"20",X"FF",X"FF",X"30",X"FF",X"30",X"60",
    X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
    X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"30",X"00",X"00",X"38",X"FF",
    X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"80",
    X"10",X"00",X"00",X"00",X"60",X"70",X"1D",X"3D",
    X"00",X"FF",X"00",X"00",X"30",X"00",X"28",X"48",
    X"30",X"00",X"28",X"38",X"00",X"00",X"00",X"30",
    X"00",X"00",X"28",X"00",X"00",X"30",X"30",X"00",
    X"10",X"00",X"FF",X"20",X"00",X"FF",X"FF",X"10",
    X"20",X"FF",X"00",X"FF",X"20",X"00",X"00",X"FF",
    X"10",X"20",X"FF",X"FF",X"00",X"00",X"FF",X"37",
    X"10",X"37",X"10",X"1D",X"18",X"00",X"00",X"00",
    X"18",X"00",X"00",X"00",X"28",X"01",X"18",X"18",
    X"01",X"28",X"01",X"30",X"10",X"FF",X"FF",X"00",
    X"00",X"00",X"18",X"00",X"00",X"00",X"70",X"80",
    X"10",X"70",X"01",X"00",X"60",X"70",X"00",X"FF",
    X"00",X"40",X"28",X"28",X"40",X"FF",X"FF",X"00",
    X"2C",X"44",X"48",X"4C",X"00",X"00",X"10",X"48",
    X"FF",X"00",X"4C",X"20",X"FF",X"24",X"00",X"18",
    X"54",X"14",X"15",X"28",X"20",X"48",X"48",X"4A",
    X"10",X"00",X"2D",X"00",X"1D",X"FF",X"FF",X"00",
    X"20",X"00",X"18",X"FF",X"10",X"20",X"FF",X"00",
    X"00",X"30",X"00",X"FF",X"37",X"10",X"37",X"10",
    X"1D",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
    X"18",X"00",X"00",X"00",X"60",X"70",X"00",X"FF",
    X"00",X"28",X"40",X"28",X"40",X"21",X"1A",X"00",
    X"00",X"00",X"FF",X"2C",X"20",X"23",X"FF",X"00",
    X"54",X"10",X"14",X"00",X"00",X"58",X"58",X"FF",
    X"00",X"5C",X"48",X"FF",X"4C",X"00",X"10",X"64",
    X"14",X"16",X"28",X"28",X"58",X"58",X"5A",X"10",
    X"10",X"14",X"00",X"00",X"00",X"10",X"10",X"00",
    X"2D",X"00",X"1D",X"FF",X"00",X"00",X"20",X"00",
    X"18",X"FF",X"10",X"20",X"FF",X"00",X"00",X"00",
    X"00",X"30",X"00",X"FF",X"37",X"10",X"37",X"10",
    X"1D",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
    X"18",X"00",X"00",X"00",X"60",X"00",X"FF",X"00",
    X"25",X"10",X"10",X"00",X"00",X"20",X"00",X"11",
    X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
    X"00",X"02",X"10",X"00",X"10",X"00",X"FF",X"18",
    X"00",X"00",X"00",X"FF",X"10",X"28",X"FF",X"00",
    X"FF",X"28",X"00",X"00",X"FF",X"10",X"28",X"FF",
    X"FF",X"00",X"FF",X"10",X"1D",X"27",X"10",X"27",
    X"10",X"00",X"00",X"00",X"10",X"FF",X"FF",X"10",
    X"00",X"00",X"00",X"02",X"00",X"60",X"70",X"00",
    X"00",X"10",X"17",X"2F",X"30",X"00",X"28",X"00",
    X"00",X"00",X"FF",X"00",X"35",X"2D",X"00",X"00",
    X"38",X"00",X"28",X"00",X"00",X"FF",X"20",X"18",
    X"00",X"20",X"28",X"28",X"00",X"00",X"10",X"00",
    X"00",X"00",X"00",X"00",X"FF",X"00",X"10",X"02",
    X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"60",
    X"70",X"00",X"10",X"00",X"10",X"60",X"70",X"00",
    X"10",X"00",X"10",X"FF",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"65",X"02",X"00",X"03",X"03",X"01",X"06",
    X"03",X"01",X"A3",X"00",X"02",X"00",X"03",X"03",
    X"01",X"05",X"03",X"01",X"A3",X"00",X"98",X"02",
    X"00",X"00",X"D3",X"B3",X"00",X"00",X"01",X"B6",
    X"70",X"01",X"03",X"60",X"70",X"01",X"06",X"03",
    X"01",X"C3",X"03",X"01",X"B3",X"03",X"03",X"01",
    X"06",X"03",X"01",X"A3",X"88",X"FF",X"C5",X"B0",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"16",X"03",X"65",X"01",
    X"00",X"05",X"B3",X"02",X"A3",X"B3",X"FF",X"A3",
    X"70",X"02",X"B3",X"B3",X"00",X"A3",X"01",X"00",
    X"05",X"70",X"02",X"B3",X"B3",X"FF",X"A3",X"00",
    X"16",X"02",X"A3",X"00",X"B3",X"01",X"A3",X"FF",
    X"02",X"05",X"00",X"00",X"00",X"16",X"02",X"B3",
    X"00",X"00",X"16",X"01",X"B3",X"80",X"05",X"88",
    X"B3",X"01",X"B3",X"00",X"16",X"80",X"98",X"A5",
    X"A6",X"00",X"00",X"70",X"01",X"B3",X"FF",X"00",
    X"05",X"20",X"02",X"00",X"03",X"01",X"A3",X"03",
    X"B3",X"01",X"05",X"03",X"01",X"C3",X"FF",X"06",
    X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",
    X"16",X"03",X"00",X"00",X"16",X"FF",X"00",X"01",
    X"00",X"03",X"00",X"03",X"00",X"70",X"FF",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"02",
    X"00",X"00",X"00",X"16",X"60",X"02",X"A3",X"00",
    X"00",X"16",X"60",X"02",X"00",X"00",X"00",X"16",
    X"60",X"01",X"A3",X"60",X"A3",X"01",X"05",X"00",
    X"16",X"01",X"03",X"03",X"01",X"B3",X"03",X"03",
    X"00",X"17",X"01",X"03",X"00",X"17",X"03",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
    X"00",X"70",X"01",X"A3",X"03",X"03",X"00",X"16",
    X"03",X"03",X"00",X"17",X"60",X"02",X"00",X"00",
    X"80",X"10",X"70",X"60",X"A0",X"01",X"90",X"05",
    X"00",X"00",X"A3",X"01",X"B3",X"20",X"02",X"05",
    X"03",X"01",X"A3",X"60",X"01",X"03",X"00",X"00",
    X"FF",X"A3",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"60",
    X"02",X"00",X"FF",X"00",X"00",X"16",X"70",X"01",
    X"00",X"03",X"03",X"00",X"16",X"03",X"03",X"00",
    X"80",X"16",X"80",X"60",X"01",X"A3",X"60",X"A3",
    X"01",X"05",X"00",X"16",X"01",X"03",X"03",X"01",
    X"B3",X"03",X"03",X"00",X"17",X"01",X"03",X"00",
    X"17",X"01",X"03",X"00",X"03",X"90",X"FF",X"00",
    X"00",X"00",X"00",X"75",X"00",X"01",X"65",X"03",
    X"03",X"70",X"B3",X"02",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
    X"02",X"A3",X"00",X"00",X"00",X"00",X"00",X"16",
    X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",
    X"16",X"00",X"00",X"00",X"03",X"01",X"00",X"FF",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"17",X"16",X"17",X"04",X"65",X"01",
    X"00",X"A3",X"E3",X"01",X"05",X"05",X"A3",X"02",
    X"C3",X"B3",X"FF",X"D3",X"00",X"17",X"17",X"04",
    X"A3",X"01",X"00",X"A3",X"C3",X"01",X"05",X"05",
    X"A3",X"02",X"D3",X"B3",X"FF",X"E3",X"16",X"A3",
    X"01",X"C3",X"07",X"A6",X"00",X"00",X"D3",X"01",
    X"A3",X"20",X"02",X"06",X"03",X"01",X"C3",X"03",
    X"D3",X"01",X"06",X"03",X"01",X"E3",X"00",X"FF",
    X"07",X"00",X"00",X"00",X"00",X"B3",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
    X"01",X"00",X"FF",X"00",X"00",X"00",X"17",X"00",
    X"00",X"00",X"17",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"B0",
    X"04",X"65",X"01",X"00",X"B3",X"E3",X"01",X"05",
    X"05",X"A3",X"02",X"C3",X"A3",X"FF",X"D3",X"00",
    X"00",X"17",X"00",X"17",X"17",X"04",X"00",X"01",
    X"00",X"B3",X"E3",X"01",X"05",X"05",X"A3",X"02",
    X"C3",X"A3",X"FF",X"D3",X"00",X"17",X"00",X"17",
    X"17",X"05",X"00",X"01",X"00",X"B3",X"E3",X"01",
    X"05",X"05",X"A3",X"02",X"C3",X"A3",X"FF",X"D3",
    X"00",X"16",X"01",X"80",X"00",X"00",X"16",X"C0",
    X"90",X"00",X"00",X"70",X"01",X"A3",X"20",X"02",
    X"05",X"03",X"01",X"A3",X"03",X"01",X"C3",X"00",
    X"FF",X"06",X"00",X"00",X"00",X"00",X"B3",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"03",X"01",X"00",X"FF",X"00",X"04",X"00",
    X"00",X"00",X"73",X"01",X"03",X"03",X"00",X"04",
    X"00",X"00",X"10",X"00",X"00",X"28",X"10",X"FF",
    X"20",X"00",X"00",X"1F",X"30",X"10",X"05",X"00",
    X"00",X"18",X"28",X"00",X"48",X"00",X"38",X"47",
    X"FF",X"10",X"FF",X"00",X"FF",X"00",X"20",X"00",
    X"FF",X"18",X"00",X"00",X"00",X"00",X"00",X"58",
    X"1F",X"30",X"10",X"05",X"00",X"00",X"18",X"28",
    X"00",X"48",X"00",X"38",X"47",X"FF",X"10",X"FF",
    X"00",X"FF",X"00",X"20",X"00",X"FF",X"18",X"00",
    X"00",X"10",X"00",X"00",X"20",X"FF",X"00",X"28",
    X"05",X"00",X"10",X"1F",X"30",X"05",X"00",X"00",
    X"18",X"28",X"00",X"48",X"00",X"38",X"FF",X"47",
    X"FF",X"00",X"FF",X"00",X"10",X"FF",X"18",X"00",
    X"00",X"10",X"1F",X"30",X"05",X"00",X"00",X"18",
    X"28",X"00",X"48",X"00",X"38",X"FF",X"47",X"FF",
    X"00",X"FF",X"00",X"10",X"FF",X"18",X"00",X"00",
    X"0F",X"0F",X"00",X"0F",X"00",X"0F",X"66",X"96",
    X"0F",X"DB",X"66",X"73",X"00",X"00",X"95",X"00",
    X"72",X"00",X"00",X"72",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal bram0 : t_bram := (
    X"01",X"00",X"00",X"08",X"00",X"04",X"00",X"08",
    X"00",X"2A",X"FD",X"04",X"AD",X"00",X"0E",X"98",
    X"10",X"14",X"18",X"1C",X"20",X"24",X"28",X"2C",
    X"30",X"34",X"38",X"3C",X"40",X"44",X"48",X"4C",
    X"50",X"54",X"00",X"FC",X"58",X"10",X"5C",X"12",
    X"60",X"00",X"20",X"00",X"10",X"00",X"24",X"90",
    X"00",X"10",X"14",X"18",X"1C",X"20",X"24",X"28",
    X"2C",X"30",X"34",X"38",X"3C",X"40",X"44",X"48",
    X"4C",X"50",X"54",X"58",X"5C",X"00",X"11",X"60",
    X"00",X"13",X"68",X"01",X"08",X"00",X"00",X"08",
    X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"3C",
    X"04",X"00",X"40",X"08",X"00",X"44",X"0C",X"00",
    X"08",X"48",X"00",X"3C",X"08",X"00",X"00",X"04",
    X"08",X"0C",X"10",X"14",X"18",X"1C",X"20",X"24",
    X"28",X"2C",X"08",X"00",X"00",X"04",X"08",X"0C",
    X"10",X"14",X"18",X"1C",X"20",X"24",X"28",X"2C",
    X"00",X"08",X"00",X"19",X"12",X"10",X"08",X"00",
    X"0C",X"08",X"00",X"FF",X"00",X"00",X"08",X"21",
    X"08",X"00",X"21",X"E8",X"00",X"0A",X"04",X"02",
    X"1B",X"0D",X"01",X"12",X"00",X"00",X"18",X"30",
    X"FF",X"00",X"12",X"00",X"00",X"02",X"1B",X"0D",
    X"12",X"ED",X"23",X"08",X"00",X"C0",X"20",X"00",
    X"00",X"05",X"02",X"1A",X"0D",X"38",X"00",X"00",
    X"08",X"04",X"3C",X"34",X"30",X"2C",X"28",X"24",
    X"1C",X"12",X"10",X"18",X"00",X"20",X"80",X"80",
    X"21",X"21",X"00",X"04",X"FD",X"00",X"27",X"21",
    X"01",X"21",X"08",X"00",X"40",X"00",X"10",X"51",
    X"0C",X"00",X"00",X"20",X"14",X"21",X"FF",X"02",
    X"80",X"21",X"00",X"FF",X"18",X"FE",X"FF",X"0C",
    X"08",X"12",X"00",X"00",X"02",X"1A",X"0D",X"10",
    X"00",X"12",X"20",X"10",X"80",X"21",X"FD",X"FE",
    X"18",X"00",X"21",X"FF",X"12",X"00",X"00",X"18",
    X"12",X"21",X"00",X"02",X"1A",X"0D",X"FE",X"10",
    X"00",X"12",X"ED",X"FC",X"23",X"FE",X"40",X"21",
    X"0C",X"08",X"10",X"02",X"1A",X"0D",X"F2",X"04",
    X"10",X"12",X"92",X"21",X"10",X"00",X"04",X"02",
    X"1A",X"0D",X"10",X"40",X"0C",X"10",X"10",X"B8",
    X"14",X"3C",X"21",X"38",X"34",X"30",X"2C",X"28",
    X"24",X"20",X"1C",X"18",X"08",X"40",X"00",X"00",
    X"26",X"00",X"08",X"00",X"00",X"00",X"C2",X"C2",
    X"7F",X"FF",X"FF",X"FF",X"24",X"80",X"24",X"2A",
    X"25",X"2E",X"25",X"23",X"1E",X"34",X"00",X"07",
    X"02",X"00",X"23",X"02",X"00",X"23",X"21",X"2C",
    X"21",X"2D",X"00",X"24",X"07",X"80",X"00",X"43",
    X"24",X"FD",X"01",X"80",X"24",X"06",X"00",X"80",
    X"40",X"24",X"FD",X"FF",X"1D",X"7F",X"FF",X"C2",
    X"24",X"C0",X"25",X"C0",X"25",X"00",X"08",X"00",
    X"23",X"1E",X"04",X"00",X"07",X"50",X"21",X"21",
    X"50",X"21",X"50",X"21",X"23",X"D5",X"00",X"00",
    X"08",X"00",X"21",X"00",X"08",X"00",X"00",X"00",
    X"26",X"00",X"3C",X"00",X"00",X"00",X"7F",X"FF",
    X"80",X"24",X"24",X"25",X"25",X"FF",X"FF",X"18",
    X"02",X"02",X"12",X"02",X"00",X"18",X"12",X"21",
    X"FF",X"18",X"02",X"12",X"FF",X"02",X"18",X"21",
    X"02",X"00",X"C2",X"12",X"21",X"21",X"21",X"40",
    X"25",X"1B",X"C2",X"FF",X"C2",X"00",X"81",X"FF",
    X"24",X"06",X"21",X"00",X"42",X"24",X"FD",X"01",
    X"0F",X"26",X"7F",X"FF",X"C2",X"24",X"C0",X"25",
    X"C0",X"25",X"00",X"08",X"00",X"00",X"08",X"00",
    X"21",X"00",X"08",X"00",X"00",X"00",X"7F",X"FF",
    X"80",X"24",X"24",X"25",X"25",X"00",X"02",X"02",
    X"1B",X"0D",X"FF",X"02",X"12",X"00",X"FF",X"18",
    X"02",X"12",X"02",X"00",X"18",X"12",X"21",X"FF",
    X"18",X"02",X"12",X"FF",X"02",X"18",X"21",X"02",
    X"00",X"02",X"12",X"21",X"21",X"21",X"00",X"25",
    X"23",X"00",X"02",X"1A",X"0D",X"12",X"21",X"1D",
    X"C2",X"FF",X"C2",X"00",X"7E",X"FF",X"24",X"06",
    X"23",X"00",X"42",X"24",X"FD",X"01",X"11",X"00",
    X"0F",X"26",X"7F",X"FF",X"C2",X"24",X"C0",X"25",
    X"C0",X"25",X"00",X"08",X"00",X"00",X"08",X"00",
    X"21",X"00",X"08",X"00",X"00",X"7F",X"FF",X"80",
    X"C2",X"24",X"25",X"FF",X"9D",X"23",X"05",X"C0",
    X"1F",X"07",X"00",X"07",X"02",X"00",X"23",X"08",
    X"00",X"44",X"21",X"20",X"21",X"21",X"00",X"24",
    X"22",X"00",X"96",X"00",X"43",X"24",X"FD",X"01",
    X"80",X"24",X"07",X"7F",X"80",X"40",X"24",X"FD",
    X"FF",X"7F",X"FF",X"24",X"C0",X"C2",X"25",X"C0",
    X"25",X"00",X"08",X"00",X"23",X"E1",X"00",X"21",
    X"00",X"08",X"00",X"58",X"96",X"00",X"00",X"00",
    X"1E",X"21",X"C2",X"C2",X"2B",X"1D",X"2B",X"19",
    X"00",X"02",X"FF",X"01",X"C2",X"C2",X"FF",X"FF",
    X"2B",X"0D",X"2B",X"11",X"7F",X"FF",X"24",X"24",
    X"80",X"25",X"25",X"2B",X"02",X"00",X"23",X"08",
    X"00",X"08",X"01",X"08",X"FF",X"08",X"23",X"75",
    X"00",X"75",X"00",X"75",X"00",X"75",X"00",X"00",
    X"00",X"00",X"26",X"08",X"2B",X"00",X"00",X"00",
    X"26",X"08",X"2B",X"B8",X"01",X"24",X"20",X"1C",
    X"18",X"14",X"44",X"40",X"34",X"30",X"2C",X"28",
    X"3C",X"06",X"4B",X"38",X"06",X"86",X"94",X"86",
    X"06",X"8E",X"86",X"00",X"4B",X"64",X"06",X"86",
    X"94",X"86",X"06",X"8E",X"86",X"00",X"21",X"DA",
    X"0A",X"00",X"06",X"86",X"1A",X"01",X"8E",X"86",
    X"00",X"94",X"06",X"00",X"00",X"8E",X"06",X"86",
    X"DC",X"06",X"86",X"8E",X"06",X"06",X"86",X"94",
    X"06",X"06",X"8E",X"86",X"21",X"E3",X"86",X"06",
    X"44",X"3C",X"34",X"2C",X"24",X"20",X"1C",X"18",
    X"14",X"40",X"38",X"30",X"28",X"08",X"48",X"C0",
    X"00",X"34",X"30",X"2C",X"28",X"24",X"20",X"1C",
    X"18",X"14",X"3C",X"38",X"E0",X"1A",X"86",X"8E",
    X"00",X"86",X"06",X"75",X"86",X"06",X"F8",X"86",
    X"00",X"75",X"06",X"06",X"0A",X"86",X"3C",X"00",
    X"86",X"00",X"75",X"06",X"06",X"F8",X"86",X"00",
    X"E4",X"75",X"86",X"43",X"06",X"8E",X"86",X"FF",
    X"4B",X"86",X"00",X"00",X"00",X"EC",X"75",X"06",
    X"07",X"00",X"E4",X"8E",X"86",X"00",X"86",X"26",
    X"06",X"94",X"86",X"00",X"E8",X"00",X"26",X"86",
    X"06",X"02",X"0C",X"00",X"94",X"06",X"FF",X"18",
    X"86",X"12",X"4B",X"02",X"86",X"94",X"06",X"86",
    X"06",X"DC",X"06",X"86",X"3C",X"06",X"EC",X"06",
    X"3C",X"34",X"2C",X"00",X"24",X"20",X"1C",X"18",
    X"14",X"38",X"30",X"28",X"06",X"94",X"40",X"00",
    X"E8",X"3D",X"00",X"00",X"EC",X"E8",X"14",X"8E",
    X"00",X"06",X"14",X"07",X"18",X"00",X"D0",X"10",
    X"1C",X"18",X"14",X"2C",X"28",X"24",X"00",X"75",
    X"20",X"63",X"00",X"E8",X"00",X"75",X"86",X"29",
    X"00",X"F8",X"00",X"75",X"00",X"2C",X"00",X"FC",
    X"00",X"8E",X"86",X"00",X"86",X"94",X"86",X"00",
    X"E8",X"3C",X"86",X"86",X"DC",X"06",X"85",X"06",
    X"00",X"00",X"3C",X"86",X"00",X"04",X"06",X"2C",
    X"24",X"1C",X"18",X"14",X"10",X"28",X"20",X"8E",
    X"30",X"00",X"DC",X"06",X"85",X"06",X"00",X"EC",
    X"B7",X"86",X"00",X"08",X"00",X"75",X"00",X"37",
    X"00",X"26",X"00",X"00",X"00",X"94",X"21",X"86",
    X"03",X"0F",X"06",X"94",X"86",X"21",X"4B",X"06",
    X"86",X"DC",X"06",X"00",X"3C",X"86",X"02",X"00",
    X"F2",X"06",X"2C",X"24",X"1C",X"00",X"18",X"14",
    X"10",X"28",X"20",X"08",X"30",X"00",X"F0",X"00",
    X"75",X"00",X"9E",X"00",X"00",X"E8",X"00",X"DC",
    X"00",X"85",X"06",X"00",X"F4",X"B7",X"86",X"00",
    X"00",X"FC",X"26",X"00",X"8E",X"86",X"00",X"86",
    X"94",X"86",X"00",X"E8",X"3C",X"86",X"86",X"DC",
    X"06",X"85",X"06",X"00",X"00",X"3C",X"86",X"00",
    X"04",X"8E",X"06",X"00",X"EA",X"26",X"D0",X"1C",
    X"2C",X"28",X"24",X"86",X"20",X"DC",X"06",X"85",
    X"06",X"00",X"06",X"75",X"10",X"10",X"08",X"00",
    X"2C",X"24",X"1C",X"28",X"20",X"08",X"30",X"00",
    X"75",X"06",X"10",X"0A",X"00",X"2C",X"24",X"E4",
    X"1C",X"28",X"20",X"06",X"3C",X"30",X"2C",X"24",
    X"E4",X"1C",X"28",X"20",X"06",X"8E",X"30",X"B8",
    X"00",X"18",X"14",X"34",X"30",X"00",X"00",X"14",
    X"00",X"44",X"40",X"3C",X"38",X"2C",X"28",X"24",
    X"20",X"1C",X"0C",X"E8",X"10",X"76",X"06",X"94",
    X"00",X"06",X"86",X"3C",X"86",X"06",X"06",X"75",
    X"86",X"06",X"F4",X"86",X"00",X"10",X"18",X"89",
    X"06",X"94",X"00",X"06",X"86",X"3C",X"86",X"06",
    X"06",X"75",X"86",X"06",X"F4",X"86",X"E8",X"86",
    X"3C",X"06",X"06",X"86",X"02",X"0F",X"06",X"94",
    X"86",X"21",X"4B",X"86",X"86",X"94",X"06",X"86",
    X"06",X"DC",X"06",X"86",X"3C",X"06",X"01",X"EE",
    X"06",X"44",X"3C",X"34",X"24",X"86",X"2C",X"1C",
    X"18",X"14",X"40",X"38",X"30",X"28",X"20",X"06",
    X"94",X"48",X"B8",X"00",X"34",X"30",X"24",X"00",
    X"3C",X"38",X"1C",X"00",X"44",X"40",X"2C",X"28",
    X"24",X"20",X"1C",X"18",X"14",X"10",X"20",X"00",
    X"D9",X"06",X"94",X"00",X"06",X"86",X"3C",X"06",
    X"86",X"06",X"75",X"86",X"06",X"F4",X"86",X"00",
    X"00",X"30",X"00",X"2C",X"28",X"EE",X"00",X"94",
    X"00",X"06",X"86",X"3C",X"06",X"86",X"06",X"75",
    X"86",X"06",X"F4",X"86",X"00",X"14",X"00",X"28",
    X"2C",X"02",X"00",X"94",X"00",X"06",X"86",X"8E",
    X"06",X"86",X"06",X"75",X"86",X"06",X"F4",X"86",
    X"00",X"E8",X"8E",X"00",X"00",X"00",X"F0",X"00",
    X"26",X"01",X"0E",X"00",X"94",X"06",X"21",X"4B",
    X"06",X"86",X"DC",X"06",X"86",X"3C",X"06",X"01",
    X"F2",X"06",X"44",X"3C",X"34",X"24",X"86",X"2C",
    X"1C",X"18",X"14",X"10",X"40",X"38",X"30",X"28",
    X"20",X"06",X"3C",X"48",X"E0",X"1C",X"BA",X"10",
    X"10",X"00",X"06",X"94",X"86",X"06",X"1C",X"57",
    X"20",X"07",X"21",X"01",X"02",X"42",X"21",X"FB",
    X"40",X"08",X"00",X"C0",X"21",X"21",X"53",X"20",
    X"11",X"25",X"42",X"02",X"2B",X"01",X"42",X"80",
    X"F7",X"40",X"F5",X"02",X"F3",X"00",X"23",X"01",
    X"F1",X"25",X"08",X"00",X"1F",X"00",X"20",X"21",
    X"C0",X"21",X"21",X"70",X"20",X"11",X"25",X"42",
    X"02",X"2B",X"01",X"42",X"80",X"F7",X"40",X"F5",
    X"02",X"F3",X"00",X"23",X"01",X"F1",X"25",X"02",
    X"00",X"23",X"08",X"00",X"23",X"E2",X"01",X"23",
    X"68",X"01",X"21",X"C0",X"21",X"92",X"20",X"0F",
    X"25",X"42",X"02",X"2B",X"01",X"42",X"F8",X"80",
    X"F6",X"02",X"F4",X"00",X"23",X"F3",X"25",X"08",
    X"00",X"21",X"C0",X"21",X"A9",X"20",X"0F",X"25",
    X"42",X"02",X"2B",X"01",X"42",X"F8",X"80",X"F6",
    X"02",X"F4",X"00",X"23",X"F3",X"25",X"08",X"00",
    X"DA",X"DA",X"00",X"DA",X"00",X"DA",X"66",X"B5",
    X"DA",X"55",X"66",X"26",X"00",X"00",X"55",X"00",
    X"18",X"00",X"00",X"18",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );

-- This is a 16-bit SRAM split in 2 byte slices; so each slice will have two
-- bytes for each word of SRAM_SIZE
type t_sram is array(0 to SRAM_SIZE*2-1) of std_logic_vector(7 downto 0);
signal sram1 : t_sram := (
    X"00",X"27",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal sram0 : t_sram := (
    X"00",X"10",X"00",X"38",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );


signal data_uart :          std_logic_vector(31 downto 0);
signal data_uart_status :   std_logic_vector(31 downto 0);
signal uart_tx_rdy :        std_logic := '1';
signal uart_rx_rdy :        std_logic := '1';

--------------------------------------------------------------------------------

signal clk :                std_logic := '0';
signal reset :              std_logic := '1';
signal interrupt :          std_logic := '0';
signal done :               std_logic := '0';

-- interface to asynchronous 16-bit-wide external SRAM
signal sram_address :       std_logic_vector(SRAM_ADDR_SIZE-1 downto 1);
signal sram_databus :       std_logic_vector(15 downto 0);
signal sram_byte_we_n :     std_logic_vector(1 downto 0);
signal sram_oe_n :          std_logic;

-- interface cpu-cache
signal cpu_data_rd_addr :   t_word;
signal cpu_data_rd_vma :    std_logic;
signal cpu_data_rd :        t_word;
signal cpu_code_rd_addr :   t_pc;
signal cpu_code_rd :        t_word;
signal cpu_code_rd_vma :    std_logic;
signal cpu_data_wr_addr :   t_pc;
signal cpu_data_wr :        t_word;
signal cpu_byte_we :        std_logic_vector(3 downto 0);
signal cpu_mem_wait :       std_logic;

-- interface to i/o
signal io_rd_data :         std_logic_vector(31 downto 0);
signal io_wr_data :         std_logic_vector(31 downto 0);
signal io_rd_addr :         std_logic_vector(31 downto 2);
signal io_wr_addr :         std_logic_vector(31 downto 2);
signal io_rd_vma :          std_logic;
signal io_byte_we :         std_logic_vector(3 downto 0);


--------------------------------------------------------------------------------
-- Logging signals

-- These are internal CPU signal mirrored using Modelsim's SignalSpy
signal rbank :              t_rbank;
signal pc, cp0_epc :        std_logic_vector(31 downto 2);
signal reg_hi, reg_lo :     t_word;
signal negate_reg_lo :      std_logic;
signal ld_upper_byte :      std_logic;
signal ld_upper_hword :     std_logic;
signal data_rd_vma :        std_logic;
signal code_rd_vma :        std_logic;
signal data_rd_address :    std_logic_vector(31 downto 0);


-- Log file
file l_file: TEXT open write_mode is "hw_sim_log.txt";

-- Console output log file
file con_file: TEXT open write_mode is "hw_sim_console_log.txt";

-- Maximum line size of for console output log. Lines longer than this will be
-- truncated.
constant CONSOLE_LOG_LINE_SIZE : integer := 1024*4;

-- Console log line buffer
signal con_line_buf :       string(1 to CONSOLE_LOG_LINE_SIZE);
signal con_line_ix :        integer := 1;

-- Debug signals ---------------------------------------------------------------


signal full_rd_addr :       std_logic_vector(31 downto 0);
signal full_wr_addr :       std_logic_vector(31 downto 0);
signal full_code_addr :     std_logic_vector(31 downto 0);


begin

    cpu: entity work.mips_cpu
    port map (
        interrupt   => '0',
        
        data_rd_addr=> cpu_data_rd_addr,
        data_rd_vma => cpu_data_rd_vma,
        data_rd     => cpu_data_rd,
        
        code_rd_addr=> cpu_code_rd_addr,
        code_rd     => cpu_code_rd,
        code_rd_vma => cpu_code_rd_vma,
        
        data_wr_addr=> cpu_data_wr_addr,
        data_wr     => cpu_data_wr,
        byte_we     => cpu_byte_we,

        mem_wait    => cpu_mem_wait,
        
        clk         => clk,
        reset       => reset
    );

    cache: entity work.mips_cache_stub
    generic map (
        BRAM_ADDR_SIZE => BRAM_ADDR_SIZE,
        SRAM_ADDR_SIZE => SRAM_ADDR_SIZE
    )
    port map (
        clk             => clk,
        reset           => reset,
        
        -- Interface to CPU core
        data_rd_addr    => cpu_data_rd_addr,
        data_rd         => cpu_data_rd,
        data_rd_vma     => cpu_data_rd_vma,
                        
        code_rd_addr    => cpu_code_rd_addr,
        code_rd         => cpu_code_rd,
        code_rd_vma     => cpu_code_rd_vma,
                        
        data_wr_addr    => cpu_data_wr_addr,
        byte_we         => cpu_byte_we,
        data_wr         => cpu_data_wr,
                        
        mem_wait        => cpu_mem_wait,
        
        -- interface to FPGA i/o devices
        io_rd_data      => io_rd_data,
        io_wr_data      => io_wr_data,
        io_rd_addr      => io_rd_addr,
        io_wr_addr      => io_wr_addr,
        io_rd_vma       => io_rd_vma,
        io_byte_we      => io_byte_we,

        -- interface to synchronous 32-bit-wide FPGA BRAM
        bram_rd_data    => bram_rd_data,
        bram_wr_data    => bram_wr_data,
        bram_rd_addr    => bram_rd_addr,
        bram_wr_addr    => bram_wr_addr,
        bram_byte_we    => bram_byte_we,
        
        -- interface to asynchronous 16-bit-wide external SRAM
        sram_address    => sram_address,
        sram_databus    => sram_databus,
        sram_byte_we_n  => sram_byte_we_n,
        sram_oe_n       => sram_oe_n
    );

    ---------------------------------------------------------------------------
    -- Master clock: free running clock used as main module clock
    run_master_clock:
    process(done, clk)
    begin
        if done = '0' then
            clk <= not clk after T/2;
        end if;
    end process run_master_clock;

    drive_uut:
    process
    variable l : line;
    begin
        wait for T*4;
        reset <= '0';
        
        wait for T*SIMULATION_LENGTH;

        -- Flush console output to log console file (in case the end of the
        -- simulation caugh an unterminated line in the buffer)
        if con_line_ix > 1 then
            write(l, con_line_buf(1 to con_line_ix));
            writeline(con_file, l);
        end if;

        print("TB0 finished");
        done <= '1';
        wait;
        
    end process drive_uut;

    full_rd_addr <= cpu_data_rd_addr;
    full_wr_addr <= cpu_data_wr_addr & "00";
    full_code_addr <= cpu_code_rd_addr & "00";

    data_ram_block:
    process(clk)
    begin
        if clk'event and clk='1' then
            if reset='0' then
                bram_rd_data <= 
                    bram3(conv_integer(unsigned(bram_rd_addr))) &
                    bram2(conv_integer(unsigned(bram_rd_addr))) &
                    bram1(conv_integer(unsigned(bram_rd_addr))) &
                    bram0(conv_integer(unsigned(bram_rd_addr)));
                
                if bram_byte_we(3)='1' then
                    bram3(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr(31 downto 24);
                end if;
                if bram_byte_we(2)='1' then
                    bram2(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr(23 downto 16);
                end if;
                if bram_byte_we(1)='1' then
                    bram1(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr(15 downto  8);
                end if;
                if bram_byte_we(0)='1' then
                    bram0(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr( 7 downto  0);
                end if;
            end if;
        end if;
    end process data_ram_block;

    sram_databus <=
        sram1(conv_integer(unsigned(sram_address))) &
        sram0(conv_integer(unsigned(sram_address)))   when sram_oe_n='0'
        else (others => 'Z');

    -- Do a very basic simulation of an external SRAM
    simulated_sram:
    process(sram_byte_we_n, sram_address)
    begin
        -- FIXME should add OE\ to control logic
        if sram_byte_we_n'event or sram_address'event then
            if sram_byte_we_n(1)='0' then
                sram1(conv_integer(unsigned(sram_address))) <= sram_databus(15 downto  8);
            end if;
            if sram_byte_we_n(0)='0' then
                sram0(conv_integer(unsigned(sram_address))) <= sram_databus( 7 downto  0);
            end if;
        end if;
    end process simulated_sram;


    simulated_io:
    process(clk)
    variable i : integer;
    variable uart_data : integer;
    begin
        if clk'event and clk='1' then
            
            if io_byte_we/="0000" then
                if io_wr_addr(31 downto 28)=X"2" then
                    -- Write to UART
                    
                    -- If we're simulating the UART TX time, pulse RDY low
                    if SIMULATED_UART_TX_TIME > 0 us then
                        uart_tx_rdy <= '0', '1' after SIMULATED_UART_TX_TIME;
                    end if;
                    
                    -- TX data may come from the high or low byte (opcodes.s
                    -- uses high byte, no_op.c uses low)
                    if io_byte_we(0)='1' then
                        uart_data := conv_integer(unsigned(io_wr_data(7 downto 0)));
                    else
                        uart_data := conv_integer(unsigned(io_wr_data(31 downto 24)));
                    end if;
                    
                    -- UART TX data goes to output after a bit of line-buffering
                    -- and editing
                    if uart_data = 10 then
                        -- CR received: print output string and clear it
                        print(con_file, con_line_buf(1 to con_line_ix));
                        con_line_ix <= 1;
                        for i in 1 to con_line_buf'high loop
                           con_line_buf(i) <= ' ';
                        end loop;
                    elsif uart_data = 13 then
                        -- ignore LF
                    else
                        -- append char to output string
                        if con_line_ix < con_line_buf'high then
                            con_line_buf(con_line_ix) <= character'val(uart_data);
                            con_line_ix <= con_line_ix + 1;
                        end if;
                    end if;
                end if;
            end if;
        end if;
    end process simulated_io;

    -- UART read registers; only status, and hardwired, for the time being
    data_uart <= data_uart_status;
    data_uart_status <= X"0000000" & "00" & uart_tx_rdy & uart_rx_rdy;


    signalspy_rbank:
    process
    begin
        init_signal_spy("/mips_tb2/cpu/p1_rbank", "rbank", 0, -1);
        init_signal_spy("/mips_tb2/cpu/p0_pc_reg", "pc", 0, -1);
        init_signal_spy("/mips_tb2/cpu/mult_div/upper_reg", "reg_hi", 0, -1);
        init_signal_spy("/mips_tb2/cpu/mult_div/lower_reg", "reg_lo", 0, -1);
        init_signal_spy("/mips_tb2/cpu/mult_div/negate_reg", "negate_reg_lo", 0, -1);
        init_signal_spy("/mips_tb2/cpu/cp0_epc", "cp0_epc", 0, -1);
        init_signal_spy("/mips_tb2/cpu/p2_ld_upper_byte", "ld_upper_byte", 0, -1);
        init_signal_spy("/mips_tb2/cpu/p2_ld_upper_byte", "ld_upper_hword", 0, -1);
        init_signal_spy("/mips_tb2/cpu/data_rd_vma", "data_rd_vma", 0, -1);
        init_signal_spy("/mips_tb2/cpu/code_rd_vma", "code_rd_vma", 0, -1);
        wait;
    end process signalspy_rbank;


    log_cpu_activity:
    process(clk)
    variable prev_rbank : t_rbank := (others => X"00000000");
    variable ri : std_logic_vector(7 downto 0);
    variable full_pc : t_word := (others => '0');
    variable prev_pc : t_word := (others => '0');
    variable prev_hi : t_word := (others => '0');
    variable prev_lo : t_word := (others => '0');
    variable prev_epc : std_logic_vector(31 downto 2) := (others => '0');
    variable wr_data : t_word := (others => '0');
    variable temp : t_word := (others => '0');
    variable size : std_logic_vector(7 downto 0) := X"00";
    variable prev_vma_data : std_logic := '0';
    variable prev_rd_addr : t_word := (others => '0');
    variable prev_rd_data : t_word := (others => '0');
    variable rd_size : std_logic_vector(7 downto 0) := X"00";
    begin
        -- we'll be sampling control & data signals at falling edge, when 
        -- they're stable
        if clk'event and clk='0' then
            if reset='0' then
                -- log loads (data only)
                -- IMPORTANT: memory reads should be logged first because we're
                -- logging them the cycle after they actually happen. If you put
                -- the log code after any other log, the order of the operations 
                -- will appear wrong in the log even though it is not.
                if prev_vma_data='1' and cpu_mem_wait='0' then
                    if ld_upper_hword='1' then
                        rd_size := X"04";
                    elsif ld_upper_byte='1' then
                        rd_size := X"02";
                    else
                        rd_size := X"01";
                    end if;
                    print(l_file, "("& hstr(prev_pc) &") ["& hstr(prev_rd_addr) &"] <"&
                          "**"&
                          --hstr(rd_size)& 
                          ">="& hstr(cpu_data_rd)& " RD");
                end if;
                
                prev_rd_data := cpu_data_rd;
                if cpu_mem_wait='0' then
                    prev_vma_data := data_rd_vma;
                    prev_rd_addr := full_rd_addr;
                end if;
                
                -- log register changes
                ri := X"00";
                for i in 0 to 31 loop
                    if prev_rbank(i)/=rbank(i) then
                        print(l_file, "("& hstr(full_pc)& ") ["& hstr(ri)& "]="& hstr(rbank(i)));
                    end if;
                    ri := ri + 1;
                end loop;

                -- log aux register changes, only when pipeline is not stalled
                if prev_lo /= reg_lo and reg_lo(0)/='U' and code_rd_vma='1' then
                    -- we're observing the value of reg_lo, but the mult core
                    -- will output the negated value in some cases. We
                    -- have to mimic that behavior.
                    if negate_reg_lo='1' then
                        -- negate reg_lo before displaying
                        prev_lo := not reg_lo;
                        prev_lo := prev_lo + 1;
                        print(l_file, "("& hstr(full_pc)& ") [LO]="& hstr(prev_lo));
                    else
                        print(l_file, "("& hstr(full_pc)& ") [LO]="& hstr(reg_lo));
                    end if;
                end if;
                if prev_hi /= reg_hi and reg_hi(0)/='U' and code_rd_vma='1' then
                    print(l_file, "("& hstr(full_pc)& ") [HI]="& hstr(reg_hi));
                end if;                
                if prev_epc /= cp0_epc and cp0_epc(31)/='U'  then
                    temp := cp0_epc & "00";
                    print(l_file, "("& hstr(full_pc)& ") [EP]="& hstr(temp));
                end if;

                -- 'remember' last value of hi and lo only when pipeline is not
                -- stalled; that's because we don't want to be tracking the
                -- changing values when mul/div is running (because the SW 
                -- simulator doesn't)
                if code_rd_vma='1' then
                    prev_hi := reg_hi;
                    prev_lo := reg_lo;
                end if;


                full_pc := pc & "00";
                prev_pc := full_pc;
                prev_rbank := rbank;
                prev_epc := cp0_epc;
                
                -- log writes
                if cpu_byte_we/="0000" then
                    wr_data := X"00000000";
                    if cpu_byte_we(3)='1' then
                        wr_data(31 downto 24) := cpu_data_wr(31 downto 24);
                    end if;
                    if cpu_byte_we(2)='1' then
                        wr_data(23 downto 16) := cpu_data_wr(23 downto 16);
                    end if;
                    if cpu_byte_we(1)='1' then
                        wr_data(15 downto  8) := cpu_data_wr(15 downto  8);
                    end if;
                    if cpu_byte_we(0)='1' then
                        wr_data( 7 downto  0) := cpu_data_wr( 7 downto  0);
                    end if;
                    size := "0000" & cpu_byte_we; -- mask, really
                    print(l_file, "("& hstr(full_pc) &") ["& hstr(full_wr_addr) &"] |"& hstr(size)& "|="& hstr(wr_data)& " WR" );
                end if;
                
                if full_code_addr(31 downto 28)="1111" then
                    print(l_file, "ERROR: Code addressed upper memory area" );
                end if;

            end if;
        end if;
    end process log_cpu_activity;
    
end architecture testbench;
