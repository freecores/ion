--##############################################################################
-- This file was generated automatically from '/src/mips_tb0_template.vhdl'.
-- 
--------------------------------------------------------------------------------
-- Simulation test bench TB0 -- not synthesizable.
--
-- Simulates the CPU core connected to a single memory block initialized with
-- the program object code and (initialized) data. The makefile for the source 
-- samples include targets to build simulation test benches using this template.
--
-- The memory setup is meant to test the 'bare' cpu, without cache and with 
-- all object code in a single 3-port memory block. 
-- Address decoding is harcoded to that of Plasma system, for the time being.
-- 
-- Console output (at addresses compatible to Plasma's) is logged to text file
-- "hw_sim_console_log.txt".
-- IMPORTANT: The code that echoes UART TX data to the simulation console does
-- line buffering; it will not print anything until it gets a CR (0x0d), and
-- will ifnore LFs (0x0a). Bear this in mind if you see no output when you 
-- expect it.
--
-- WARNING: Will only work on Modelsim; uses custom library SignalSpy.
--##############################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use std.textio.all;

use work.mips_pkg.all;
use work.mips_tb_pkg.all;
use work.txt_util.all;


entity mips_tb1 is
end mips_tb1;

architecture testbench of mips_tb1 is

--------------------------------------------------------------------------------
-- Simulation parameters

-- Master clock period
constant T : time           := 20 ns;
-- Time the UART is unavailable after writing to the TX register
-- WARNING: slite does not simulate this. The logs may be different when > 0.0!
constant SIMULATED_UART_TX_TIME : time := 0.0 us;

-- Simulation length in clock cycles 
-- 2000 is enough for 'hello' sample, 22000 enough for 10 digits of pi
constant SIMULATION_LENGTH : integer := 3000;

               
--------------------------------------------------------------------------------
-- UUT & interface signals

signal rd_addr :            std_logic_vector(31 downto 0);
signal prev_rd_addr :       std_logic_vector(31 downto 0);
signal vma_data :           std_logic;
signal vma_code :           std_logic;
signal wr_addr :            std_logic_vector(31 downto 2);
signal full_rd_addr :       std_logic_vector(31 downto 0);
signal full_wr_addr :       std_logic_vector(31 downto 0);
signal byte_we :            std_logic_vector(3 downto 0);
signal data_r :             std_logic_vector(31 downto 0);
signal data_ram :           std_logic_vector(31 downto 0);
signal data_uart :          std_logic_vector(31 downto 0);
signal data_uart_status :   std_logic_vector(31 downto 0);
signal uart_tx_rdy :        std_logic := '1';
signal uart_rx_rdy :        std_logic := '1';
signal data_w :             std_logic_vector(31 downto 0);
signal mem_wait :           std_logic := '0';
signal interrupt :          std_logic := '0';
signal code_addr :          std_logic_vector(31 downto 2);
signal full_code_addr :     std_logic_vector(31 downto 0);
signal code_r :             std_logic_vector(31 downto 0);

--------------------------------------------------------------------------------

signal clk :                std_logic := '0';
signal reset :              std_logic := '1';
signal done :               std_logic := '0';
signal test :               integer := 0;

--------------------------------------------------------------------------------
-- Logging signals

-- These are internal CPU signal mirrored using Modelsim's SignalSpy
--signal rbank :              t_rbank;
--signal pc, cp0_epc :        std_logic_vector(31 downto 2);
--signal reg_hi, reg_lo :     t_word;
--signal negate_reg_lo :      std_logic;
--signal ld_upper_byte :      std_logic;
--signal ld_upper_hword :     std_logic;
  
signal log_info :           t_log_info;  
  
-- Log file
file log_file: TEXT open write_mode is "hw_sim_log.txt";

-- Console output log file
file con_file: TEXT open write_mode is "hw_sim_console_log.txt";

-- Maximum line size of for console output log. Lines longer than this will be
-- truncated.
constant CONSOLE_LOG_LINE_SIZE : integer := 1024*4;

-- Console log line buffer
signal con_line_buf :       string(1 to CONSOLE_LOG_LINE_SIZE);
signal con_line_ix :        integer := 1;


--------------------------------------------------------------------------------

constant MEM_SIZE : integer := 1024;
constant ADDR_SIZE : integer := 10;

subtype t_address is std_logic_vector(ADDR_SIZE-1 downto 0);

signal addr_rd, addr_wr :   t_address;
signal addr_code :          t_address;

type t_code_ram is array(0 to MEM_SIZE-1) of std_logic_vector(7 downto 0);

subtype t_data_address is std_logic_vector(ADDR_SIZE-1 downto 0);
signal data_addr_rd :       t_data_address; 
signal data_addr_wr :       t_data_address;
signal code_addr_rd :       t_data_address;


-- ram0 is LSB, ram3 is MSB
signal ram3 : t_code_ram := (
    X"3C",X"27",X"3C",X"24",X"3C",X"24",X"00",X"00",
    X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
    X"33",X"34",X"13",X"23",X"13",X"23",X"17",X"00",
    X"08",X"20",X"08",X"20",X"08",X"20",X"08",X"20",
    X"40",X"40",X"00",X"33",X"17",X"23",X"03",X"00",
    X"23",X"03",X"24",X"24",X"00",X"00",X"00",X"40",
    X"3C",X"34",X"34",X"34",X"34",X"A2",X"A2",X"A2",
    X"A2",X"A2",X"A2",X"A2",X"A2",X"34",X"A2",X"34",
    X"A2",X"34",X"A2",X"34",X"A2",X"34",X"A2",X"A2",
    X"A2",X"34",X"A2",X"34",X"34",X"00",X"A2",X"A2",
    X"A2",X"34",X"A2",X"34",X"20",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"24",X"A2",X"A2",X"A2",X"34",
    X"A2",X"34",X"34",X"00",X"A2",X"A2",X"A2",X"34",
    X"A2",X"34",X"34",X"14",X"00",X"00",X"24",X"14",
    X"3C",X"14",X"00",X"00",X"00",X"00",X"00",X"A2",
    X"00",X"20",X"A2",X"24",X"34",X"14",X"00",X"00",
    X"24",X"14",X"3C",X"14",X"00",X"00",X"00",X"00",
    X"00",X"00",X"A2",X"34",X"24",X"14",X"00",X"00",
    X"24",X"14",X"3C",X"14",X"00",X"00",X"00",X"00",
    X"00",X"00",X"A2",X"24",X"24",X"14",X"00",X"00",
    X"24",X"14",X"3C",X"14",X"00",X"00",X"00",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"34",X"14",
    X"00",X"00",X"00",X"00",X"00",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"34",X"00",X"00",X"00",X"A2",
    X"24",X"34",X"00",X"00",X"00",X"00",X"00",X"20",
    X"A2",X"34",X"24",X"00",X"00",X"00",X"00",X"00",
    X"20",X"A2",X"24",X"24",X"00",X"00",X"00",X"00",
    X"20",X"A2",X"3C",X"34",X"3C",X"34",X"00",X"00",
    X"24",X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"34",
    X"00",X"00",X"00",X"A2",X"A2",X"A2",X"34",X"A2",
    X"34",X"34",X"00",X"20",X"A2",X"00",X"20",X"A2",
    X"24",X"00",X"20",X"A2",X"00",X"20",X"A2",X"24",
    X"00",X"20",X"A2",X"00",X"20",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"28",X"20",X"A2",X"28",X"20",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"2C",X"20",
    X"A2",X"2C",X"20",X"A2",X"A2",X"A2",X"34",X"A2",
    X"34",X"34",X"00",X"20",X"A2",X"00",X"20",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"34",X"00",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"34",X"00",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"A2",X"34",X"A2",
    X"34",X"A2",X"34",X"A2",X"34",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"34",X"10",X"A2",X"A2",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"34",X"34",X"34",
    X"34",X"34",X"04",X"A2",X"A2",X"10",X"A2",X"A2",
    X"A2",X"03",X"A2",X"A2",X"A2",X"A2",X"34",X"A2",
    X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"10",
    X"A2",X"A2",X"10",X"A2",X"A2",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"34",X"34",X"34",X"34",X"34",
    X"3C",X"34",X"34",X"04",X"A2",X"A2",X"04",X"A2",
    X"A2",X"04",X"00",X"A2",X"A2",X"A2",X"A2",X"34",
    X"A2",X"34",X"34",X"34",X"34",X"34",X"34",X"3C",
    X"34",X"04",X"00",X"A2",X"04",X"00",X"A2",X"10",
    X"A2",X"A2",X"A2",X"03",X"A2",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"34",X"34",X"34",X"34",X"3C",
    X"34",X"1C",X"A2",X"A2",X"1C",X"A2",X"A2",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"34",X"34",X"34",
    X"34",X"3C",X"34",X"18",X"A2",X"A2",X"18",X"A2",
    X"A2",X"18",X"00",X"A2",X"A2",X"A2",X"A2",X"34",
    X"A2",X"34",X"34",X"34",X"34",X"34",X"34",X"3C",
    X"34",X"34",X"04",X"A2",X"A2",X"04",X"A2",X"A2",
    X"04",X"00",X"A2",X"A2",X"A2",X"A2",X"34",X"A2",
    X"34",X"34",X"34",X"34",X"34",X"34",X"3C",X"34",
    X"04",X"00",X"A2",X"04",X"00",X"A2",X"10",X"A2",
    X"A2",X"A2",X"03",X"A2",X"A2",X"A2",X"A2",X"34",
    X"A2",X"34",X"34",X"34",X"34",X"34",X"34",X"34",
    X"14",X"A2",X"A2",X"14",X"A2",X"A2",X"A2",X"A2",
    X"A2",X"34",X"A2",X"34",X"34",X"34",X"08",X"A2",
    X"A2",X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"34",
    X"34",X"34",X"34",X"34",X"0C",X"A2",X"A2",X"10",
    X"A2",X"A2",X"A2",X"03",X"A2",X"A2",X"A2",X"A2",
    X"34",X"A2",X"34",X"34",X"34",X"34",X"34",X"34",
    X"3C",X"24",X"00",X"A2",X"A2",X"10",X"A2",X"A2",
    X"A2",X"03",X"A2",X"A2",X"A2",X"A2",X"34",X"A2",
    X"34",X"34",X"34",X"3C",X"24",X"00",X"A2",X"A2",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"00",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"34",X"00",X"20",
    X"A2",X"00",X"80",X"00",X"08",X"20",X"20",X"00",
    X"A2",X"08",X"00",X"00",X"08",X"00",X"20",X"A2",
    X"A2",X"34",X"A2",X"34",X"00",X"20",X"A2",X"00",
    X"80",X"00",X"08",X"20",X"20",X"00",X"08",X"00",
    X"20",X"A2",X"A2",X"34",X"A2",X"34",X"A2",X"34",
    X"A2",X"34",X"A2",X"A2",X"A2",X"34",X"A2",X"00",
    X"3C",X"34",X"AC",X"80",X"A2",X"80",X"00",X"A2",
    X"80",X"00",X"A2",X"80",X"00",X"00",X"20",X"A2",
    X"20",X"A2",X"A2",X"A2",X"34",X"A2",X"00",X"3C",
    X"34",X"AC",X"80",X"A2",X"80",X"A2",X"80",X"A2",
    X"80",X"A2",X"A2",X"A2",X"34",X"A2",X"00",X"3C",
    X"34",X"AC",X"84",X"A2",X"84",X"A2",X"A2",X"A2",
    X"34",X"A2",X"00",X"3C",X"34",X"AC",X"84",X"A2",
    X"84",X"A2",X"A2",X"A2",X"34",X"A2",X"00",X"24",
    X"AC",X"34",X"8C",X"A2",X"A2",X"A2",X"34",X"A2",
    X"34",X"A2",X"A2",X"A2",X"34",X"A2",X"00",X"34",
    X"A4",X"80",X"A2",X"80",X"A2",X"A2",X"A2",X"34",
    X"A2",X"00",X"3C",X"34",X"AC",X"80",X"A2",X"80",
    X"A2",X"80",X"A2",X"80",X"A2",X"A2",X"A2",X"34",
    X"A2",X"34",X"A2",X"34",X"A2",X"34",X"A2",X"34",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"34",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"30",X"A2",
    X"A2",X"A2",X"34",X"A2",X"3C",X"00",X"A2",X"A2",
    X"A2",X"34",X"A2",X"3C",X"34",X"3C",X"34",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"34",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"34",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"34",X"00",X"A2",
    X"A2",X"A2",X"34",X"A2",X"34",X"38",X"A2",X"A2",
    X"A2",X"34",X"A2",X"34",X"A2",X"34",X"A2",X"34",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"00",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"00",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"00",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"00",X"00",
    X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"A2",X"34",
    X"A2",X"34",X"A2",X"34",X"A2",X"A2",X"A2",X"34",
    X"A2",X"3C",X"34",X"00",X"00",X"A2",X"A2",X"A2",
    X"34",X"A2",X"3C",X"34",X"34",X"00",X"00",X"A2",
    X"A2",X"A2",X"34",X"A2",X"3C",X"34",X"00",X"A2",
    X"3C",X"00",X"20",X"A2",X"A2",X"A2",X"34",X"A2",
    X"3C",X"34",X"34",X"00",X"A2",X"34",X"3C",X"00",
    X"20",X"A2",X"A2",X"A2",X"34",X"A2",X"3C",X"34",
    X"00",X"A2",X"3C",X"00",X"A2",X"A2",X"A2",X"34",
    X"A2",X"3C",X"34",X"34",X"00",X"A2",X"34",X"3C",
    X"00",X"A2",X"A2",X"A2",X"34",X"A2",X"34",X"A2",
    X"34",X"A2",X"34",X"A2",X"A2",X"A2",X"08",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal ram2 : t_code_ram := (
    X"1C",X"9C",X"04",X"84",X"05",X"A5",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",
    X"5A",X"1B",X"5B",X"7B",X"5B",X"7B",X"5B",X"00",
    X"00",X"84",X"00",X"84",X"00",X"84",X"00",X"84",
    X"1B",X"1A",X"1A",X"5A",X"40",X"7B",X"60",X"00",
    X"7B",X"60",X"02",X"03",X"43",X"00",X"00",X"80",
    X"14",X"15",X"16",X"17",X"18",X"97",X"95",X"97",
    X"95",X"97",X"95",X"97",X"95",X"02",X"82",X"02",
    X"82",X"02",X"82",X"02",X"82",X"02",X"82",X"97",
    X"95",X"02",X"82",X"03",X"04",X"64",X"82",X"97",
    X"95",X"02",X"82",X"04",X"82",X"82",X"97",X"95",
    X"02",X"82",X"04",X"85",X"85",X"97",X"95",X"02",
    X"82",X"03",X"04",X"64",X"82",X"97",X"95",X"02",
    X"82",X"02",X"03",X"60",X"43",X"07",X"01",X"61",
    X"01",X"41",X"00",X"06",X"00",X"00",X"00",X"84",
    X"00",X"84",X"84",X"02",X"03",X"60",X"43",X"07",
    X"01",X"61",X"01",X"41",X"00",X"06",X"00",X"00",
    X"00",X"04",X"84",X"02",X"03",X"60",X"43",X"07",
    X"01",X"61",X"01",X"41",X"00",X"06",X"00",X"00",
    X"00",X"04",X"84",X"02",X"03",X"60",X"43",X"07",
    X"01",X"61",X"01",X"41",X"00",X"06",X"00",X"00",
    X"84",X"97",X"95",X"02",X"82",X"02",X"03",X"60",
    X"43",X"07",X"00",X"00",X"00",X"84",X"97",X"95",
    X"02",X"82",X"02",X"03",X"43",X"00",X"00",X"84",
    X"02",X"03",X"43",X"00",X"00",X"04",X"85",X"84",
    X"84",X"02",X"03",X"43",X"00",X"00",X"04",X"85",
    X"84",X"84",X"02",X"03",X"43",X"00",X"00",X"85",
    X"84",X"84",X"04",X"84",X"05",X"A5",X"85",X"00",
    X"C7",X"87",X"97",X"95",X"02",X"82",X"02",X"03",
    X"43",X"00",X"00",X"84",X"97",X"95",X"02",X"82",
    X"02",X"03",X"43",X"85",X"85",X"62",X"85",X"85",
    X"02",X"43",X"85",X"85",X"62",X"85",X"85",X"03",
    X"43",X"85",X"85",X"62",X"85",X"85",X"97",X"95",
    X"02",X"82",X"02",X"44",X"85",X"85",X"44",X"85",
    X"85",X"97",X"95",X"02",X"82",X"02",X"44",X"85",
    X"85",X"44",X"85",X"85",X"97",X"95",X"02",X"82",
    X"02",X"03",X"43",X"85",X"85",X"62",X"85",X"85",
    X"97",X"95",X"02",X"82",X"03",X"04",X"64",X"82",
    X"97",X"95",X"02",X"82",X"03",X"04",X"64",X"82",
    X"97",X"95",X"02",X"82",X"02",X"82",X"02",X"82",
    X"02",X"82",X"02",X"82",X"02",X"82",X"97",X"95",
    X"02",X"82",X"0A",X"0B",X"00",X"8A",X"96",X"8B",
    X"97",X"95",X"02",X"82",X"0A",X"0B",X"0C",X"0D",
    X"0E",X"0F",X"11",X"8A",X"8D",X"00",X"8E",X"8F",
    X"8B",X"E0",X"8C",X"96",X"97",X"95",X"02",X"82",
    X"0A",X"0B",X"0C",X"0D",X"02",X"03",X"04",X"43",
    X"8A",X"8B",X"64",X"8C",X"96",X"8D",X"97",X"95",
    X"02",X"82",X"0A",X"0B",X"0C",X"0D",X"0F",X"02",
    X"03",X"63",X"04",X"61",X"8A",X"8B",X"41",X"8C",
    X"96",X"01",X"00",X"8F",X"8D",X"97",X"95",X"02",
    X"82",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"03",
    X"63",X"71",X"00",X"8A",X"11",X"00",X"8D",X"00",
    X"8E",X"8F",X"8B",X"E0",X"8C",X"96",X"97",X"95",
    X"02",X"82",X"0A",X"0B",X"0C",X"0D",X"02",X"03",
    X"63",X"60",X"8A",X"8B",X"40",X"8C",X"96",X"8D",
    X"97",X"95",X"02",X"82",X"0A",X"0B",X"0C",X"0D",
    X"02",X"03",X"63",X"40",X"8A",X"8B",X"60",X"8C",
    X"96",X"00",X"00",X"96",X"8D",X"97",X"95",X"02",
    X"82",X"0A",X"0B",X"0C",X"0D",X"0E",X"02",X"03",
    X"63",X"04",X"40",X"8A",X"8B",X"60",X"8C",X"96",
    X"80",X"00",X"8D",X"8E",X"97",X"95",X"02",X"82",
    X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"03",X"63",
    X"10",X"00",X"8A",X"70",X"00",X"8D",X"00",X"8E",
    X"8F",X"8B",X"E0",X"8C",X"96",X"97",X"95",X"02",
    X"82",X"0A",X"0B",X"0C",X"0D",X"02",X"03",X"04",
    X"64",X"8A",X"8B",X"43",X"8C",X"96",X"8D",X"97",
    X"95",X"02",X"82",X"0A",X"0B",X"0F",X"00",X"8A",
    X"8F",X"8B",X"97",X"95",X"02",X"82",X"0A",X"0B",
    X"0C",X"0D",X"0E",X"0F",X"00",X"8A",X"8D",X"00",
    X"8E",X"8F",X"8B",X"E0",X"8C",X"96",X"97",X"95",
    X"02",X"82",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",
    X"03",X"63",X"60",X"8A",X"8D",X"00",X"8E",X"8F",
    X"8B",X"E0",X"8C",X"96",X"97",X"95",X"02",X"82",
    X"0A",X"0B",X"0F",X"03",X"63",X"60",X"8A",X"8F",
    X"8B",X"97",X"95",X"02",X"82",X"02",X"00",X"82",
    X"97",X"95",X"02",X"82",X"02",X"04",X"00",X"84",
    X"84",X"00",X"42",X"00",X"00",X"84",X"84",X"00",
    X"84",X"00",X"00",X"00",X"00",X"00",X"84",X"97",
    X"95",X"02",X"82",X"04",X"00",X"84",X"84",X"00",
    X"42",X"00",X"00",X"84",X"84",X"00",X"00",X"00",
    X"84",X"97",X"95",X"02",X"82",X"02",X"82",X"02",
    X"82",X"02",X"82",X"97",X"95",X"02",X"82",X"18",
    X"03",X"63",X"43",X"44",X"84",X"44",X"00",X"84",
    X"44",X"00",X"84",X"42",X"00",X"02",X"63",X"83",
    X"42",X"82",X"97",X"95",X"02",X"82",X"18",X"03",
    X"63",X"43",X"44",X"84",X"44",X"84",X"44",X"84",
    X"42",X"82",X"97",X"95",X"02",X"82",X"18",X"03",
    X"63",X"43",X"44",X"84",X"42",X"82",X"97",X"95",
    X"02",X"82",X"18",X"03",X"63",X"43",X"44",X"84",
    X"42",X"82",X"97",X"95",X"02",X"82",X"18",X"03",
    X"43",X"03",X"42",X"82",X"97",X"95",X"02",X"82",
    X"02",X"82",X"97",X"95",X"02",X"82",X"18",X"02",
    X"82",X"83",X"83",X"82",X"82",X"97",X"95",X"02",
    X"82",X"18",X"03",X"63",X"43",X"44",X"84",X"44",
    X"84",X"44",X"84",X"42",X"82",X"97",X"95",X"02",
    X"82",X"02",X"82",X"02",X"82",X"02",X"82",X"02",
    X"82",X"97",X"95",X"02",X"82",X"02",X"03",X"43",
    X"84",X"97",X"95",X"02",X"82",X"02",X"44",X"84",
    X"97",X"95",X"02",X"82",X"02",X"02",X"83",X"97",
    X"95",X"02",X"82",X"02",X"42",X"03",X"63",X"43",
    X"84",X"97",X"95",X"02",X"82",X"02",X"03",X"43",
    X"84",X"97",X"95",X"02",X"82",X"02",X"44",X"84",
    X"97",X"95",X"02",X"82",X"02",X"03",X"43",X"84",
    X"97",X"95",X"02",X"82",X"02",X"44",X"84",X"97",
    X"95",X"02",X"82",X"02",X"82",X"02",X"82",X"02",
    X"82",X"97",X"95",X"02",X"82",X"02",X"40",X"00",
    X"83",X"97",X"95",X"02",X"82",X"02",X"40",X"00",
    X"83",X"97",X"95",X"02",X"82",X"02",X"40",X"00",
    X"83",X"97",X"95",X"02",X"82",X"02",X"40",X"00",
    X"83",X"97",X"95",X"02",X"82",X"02",X"82",X"02",
    X"82",X"02",X"82",X"02",X"82",X"97",X"95",X"02",
    X"82",X"02",X"42",X"02",X"03",X"83",X"97",X"95",
    X"02",X"82",X"02",X"42",X"03",X"62",X"03",X"83",
    X"97",X"95",X"02",X"82",X"02",X"42",X"02",X"83",
    X"02",X"02",X"63",X"83",X"97",X"95",X"02",X"82",
    X"02",X"42",X"03",X"62",X"83",X"03",X"02",X"62",
    X"63",X"83",X"97",X"95",X"02",X"82",X"02",X"42",
    X"02",X"83",X"02",X"02",X"83",X"97",X"95",X"02",
    X"82",X"02",X"42",X"03",X"62",X"84",X"03",X"02",
    X"62",X"83",X"97",X"95",X"02",X"82",X"02",X"82",
    X"02",X"82",X"02",X"82",X"97",X"95",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal ram1 : t_code_ram := (
    X"00",X"8F",X"00",X"0F",X"00",X"0F",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"68",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"70",X"68",X"D7",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
    X"20",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
    X"00",X"1D",X"00",X"00",X"00",X"00",X"FF",X"00",
    X"80",X"00",X"00",X"00",X"10",X"00",X"20",X"00",
    X"20",X"00",X"00",X"FB",X"00",X"00",X"00",X"00",
    X"FF",X"00",X"80",X"00",X"00",X"00",X"10",X"00",
    X"20",X"20",X"00",X"06",X"FF",X"00",X"00",X"00",
    X"FF",X"00",X"80",X"00",X"00",X"00",X"10",X"00",
    X"20",X"20",X"00",X"FC",X"FF",X"00",X"00",X"00",
    X"FF",X"00",X"80",X"00",X"00",X"00",X"10",X"20",
    X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
    X"00",X"00",X"10",X"00",X"20",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
    X"FF",X"00",X"00",X"28",X"20",X"20",X"20",X"00",
    X"00",X"00",X"FF",X"00",X"28",X"20",X"20",X"20",
    X"00",X"00",X"FF",X"FF",X"00",X"28",X"20",X"20",
    X"00",X"00",X"FE",X"62",X"00",X"8D",X"00",X"30",
    X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",
    X"FF",X"20",X"00",X"00",X"20",X"00",X"00",X"FF",
    X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"FF",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
    X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
    X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"FF",X"12",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
    X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"12",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"09",X"F8",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
    X"00",X"02",X"00",X"00",X"02",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
    X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
    X"41",X"43",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"1A",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"41",
    X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"41",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"10",X"41",X"43",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"07",X"60",X"20",
    X"00",X"00",X"00",X"00",X"00",X"07",X"60",X"00",
    X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",
    X"00",X"00",X"00",X"F0",X"F0",X"0F",X"0F",X"20",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"F0",X"F0",X"20",X"00",
    X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"40",X"42",X"1A",X"1E",X"00",X"00",X"00",
    X"00",X"00",X"40",X"42",X"00",X"18",X"1E",X"00",
    X"00",X"00",X"00",X"00",X"40",X"42",X"1C",X"00",
    X"84",X"1E",X"FF",X"00",X"00",X"00",X"00",X"00",
    X"40",X"42",X"00",X"18",X"00",X"00",X"84",X"18",
    X"FF",X"00",X"00",X"00",X"00",X"00",X"40",X"42",
    X"1C",X"00",X"84",X"1E",X"00",X"00",X"00",X"00",
    X"00",X"40",X"42",X"00",X"20",X"00",X"00",X"84",
    X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal ram0 : t_code_ram := (
    X"01",X"10",X"00",X"20",X"00",X"20",X"00",X"00",
    X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"1F",X"08",X"09",X"01",X"05",X"01",X"07",X"00",
    X"20",X"04",X"20",X"05",X"20",X"06",X"20",X"0F",
    X"00",X"00",X"C2",X"01",X"03",X"04",X"08",X"00",
    X"04",X"08",X"03",X"04",X"18",X"00",X"00",X"00",
    X"00",X"0A",X"58",X"0D",X"80",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"41",X"00",X"72",
    X"00",X"69",X"00",X"74",X"00",X"68",X"00",X"00",
    X"00",X"61",X"00",X"05",X"3C",X"20",X"00",X"00",
    X"00",X"62",X"00",X"3C",X"05",X"00",X"00",X"00",
    X"63",X"00",X"32",X"0F",X"00",X"00",X"00",X"64",
    X"00",X"05",X"3C",X"20",X"00",X"00",X"00",X"65",
    X"00",X"DE",X"75",X"02",X"1A",X"0D",X"FF",X"04",
    X"00",X"02",X"00",X"0D",X"12",X"00",X"12",X"00",
    X"10",X"19",X"00",X"07",X"13",X"02",X"1A",X"0D",
    X"FF",X"04",X"00",X"02",X"00",X"0D",X"12",X"00",
    X"12",X"22",X"00",X"1C",X"E9",X"02",X"1A",X"0D",
    X"FF",X"04",X"00",X"02",X"00",X"0D",X"12",X"00",
    X"12",X"22",X"00",X"7F",X"F3",X"02",X"1A",X"0D",
    X"FF",X"04",X"00",X"02",X"00",X"0D",X"12",X"12",
    X"00",X"00",X"00",X"66",X"00",X"4D",X"0D",X"02",
    X"1B",X"0D",X"12",X"00",X"12",X"00",X"00",X"00",
    X"67",X"00",X"05",X"0D",X"18",X"00",X"12",X"00",
    X"FB",X"0D",X"18",X"10",X"12",X"22",X"21",X"02",
    X"00",X"05",X"F3",X"18",X"10",X"12",X"22",X"21",
    X"03",X"00",X"FB",X"F3",X"18",X"10",X"12",X"21",
    X"03",X"00",X"98",X"E5",X"06",X"B8",X"18",X"10",
    X"7A",X"00",X"00",X"00",X"68",X"00",X"05",X"0D",
    X"19",X"00",X"12",X"00",X"00",X"00",X"69",X"00",
    X"0A",X"0C",X"2A",X"40",X"00",X"2A",X"42",X"00",
    X"F0",X"2A",X"42",X"00",X"2A",X"44",X"00",X"FF",
    X"2A",X"44",X"00",X"2A",X"46",X"00",X"00",X"00",
    X"6A",X"00",X"0A",X"0C",X"40",X"00",X"08",X"42",
    X"00",X"00",X"00",X"6B",X"00",X"0A",X"0C",X"40",
    X"00",X"08",X"42",X"00",X"00",X"00",X"6C",X"00",
    X"0A",X"0C",X"2A",X"40",X"00",X"2A",X"42",X"00",
    X"00",X"00",X"6D",X"00",X"46",X"05",X"22",X"00",
    X"00",X"00",X"6E",X"00",X"46",X"05",X"22",X"00",
    X"00",X"00",X"42",X"00",X"72",X"00",X"61",X"00",
    X"6E",X"00",X"63",X"00",X"68",X"00",X"00",X"00",
    X"61",X"00",X"41",X"42",X"02",X"00",X"00",X"00",
    X"00",X"00",X"62",X"00",X"41",X"42",X"43",X"44",
    X"45",X"58",X"05",X"00",X"00",X"06",X"00",X"00",
    X"00",X"08",X"00",X"00",X"00",X"00",X"63",X"00",
    X"41",X"42",X"43",X"44",X"64",X"7B",X"7B",X"05",
    X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
    X"64",X"00",X"41",X"42",X"43",X"44",X"58",X"64",
    X"FF",X"34",X"7B",X"05",X"00",X"00",X"02",X"00",
    X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"65",
    X"00",X"41",X"42",X"43",X"44",X"45",X"58",X"FF",
    X"34",X"08",X"00",X"00",X"05",X"00",X"00",X"06",
    X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
    X"66",X"00",X"41",X"42",X"43",X"44",X"64",X"FF",
    X"34",X"05",X"00",X"00",X"02",X"00",X"00",X"00",
    X"00",X"00",X"67",X"00",X"41",X"42",X"43",X"44",
    X"64",X"FF",X"34",X"05",X"00",X"00",X"02",X"00",
    X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"68",
    X"00",X"41",X"42",X"43",X"44",X"45",X"64",X"FF",
    X"34",X"00",X"05",X"00",X"00",X"02",X"00",X"00",
    X"02",X"00",X"00",X"00",X"00",X"00",X"69",X"00",
    X"41",X"42",X"43",X"44",X"45",X"58",X"FF",X"34",
    X"08",X"00",X"00",X"05",X"00",X"00",X"06",X"00",
    X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"6A",
    X"00",X"41",X"42",X"43",X"44",X"64",X"7B",X"7B",
    X"05",X"00",X"00",X"02",X"00",X"00",X"00",X"00",
    X"00",X"6B",X"00",X"41",X"42",X"58",X"19",X"00",
    X"00",X"00",X"00",X"00",X"6C",X"00",X"41",X"42",
    X"43",X"44",X"45",X"58",X"2A",X"00",X"00",X"06",
    X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
    X"6D",X"00",X"41",X"42",X"43",X"44",X"45",X"58",
    X"00",X"00",X"09",X"00",X"00",X"06",X"00",X"00",
    X"00",X"08",X"00",X"00",X"00",X"00",X"6E",X"00",
    X"41",X"42",X"58",X"00",X"40",X"08",X"00",X"00",
    X"00",X"00",X"00",X"6F",X"00",X"41",X"00",X"00",
    X"00",X"00",X"70",X"00",X"7A",X"3B",X"0D",X"01",
    X"00",X"0D",X"10",X"0D",X"66",X"05",X"01",X"0D",
    X"00",X"6E",X"0D",X"00",X"6F",X"00",X"01",X"00",
    X"00",X"71",X"00",X"3D",X"0C",X"FF",X"00",X"0C",
    X"10",X"0C",X"7C",X"05",X"01",X"00",X"81",X"00",
    X"01",X"00",X"00",X"4C",X"00",X"6F",X"00",X"61",
    X"00",X"64",X"00",X"00",X"00",X"61",X"00",X"25",
    X"42",X"FC",X"10",X"10",X"00",X"11",X"00",X"00",
    X"12",X"00",X"00",X"13",X"00",X"03",X"45",X"00",
    X"49",X"00",X"00",X"00",X"62",X"00",X"25",X"42",
    X"44",X"10",X"10",X"00",X"11",X"00",X"12",X"00",
    X"13",X"00",X"00",X"00",X"63",X"00",X"25",X"41",
    X"42",X"10",X"10",X"00",X"12",X"00",X"00",X"00",
    X"64",X"00",X"25",X"41",X"42",X"10",X"10",X"00",
    X"12",X"00",X"00",X"00",X"65",X"00",X"25",X"41",
    X"10",X"00",X"10",X"00",X"00",X"00",X"67",X"00",
    X"41",X"00",X"00",X"00",X"68",X"00",X"25",X"42",
    X"10",X"10",X"00",X"11",X"00",X"00",X"00",X"69",
    X"00",X"25",X"42",X"44",X"10",X"10",X"00",X"11",
    X"00",X"12",X"00",X"13",X"00",X"00",X"00",X"4C",
    X"00",X"6F",X"00",X"67",X"00",X"69",X"00",X"63",
    X"00",X"00",X"00",X"61",X"00",X"41",X"F3",X"24",
    X"00",X"00",X"00",X"62",X"00",X"41",X"F3",X"00",
    X"00",X"00",X"63",X"00",X"41",X"02",X"00",X"00",
    X"00",X"64",X"00",X"FF",X"8E",X"0F",X"30",X"27",
    X"00",X"00",X"00",X"65",X"00",X"40",X"01",X"25",
    X"00",X"00",X"00",X"66",X"00",X"40",X"01",X"00",
    X"00",X"00",X"67",X"00",X"43",X"02",X"26",X"00",
    X"00",X"00",X"68",X"00",X"43",X"02",X"00",X"00",
    X"00",X"4D",X"00",X"6F",X"00",X"76",X"00",X"65",
    X"00",X"00",X"00",X"61",X"00",X"41",X"11",X"10",
    X"00",X"00",X"00",X"62",X"00",X"41",X"13",X"12",
    X"00",X"00",X"00",X"63",X"00",X"41",X"11",X"10",
    X"00",X"00",X"00",X"64",X"00",X"41",X"13",X"12",
    X"00",X"00",X"00",X"53",X"00",X"68",X"00",X"69",
    X"00",X"66",X"00",X"74",X"00",X"00",X"00",X"61",
    X"00",X"41",X"43",X"00",X"02",X"00",X"00",X"00",
    X"62",X"00",X"41",X"43",X"08",X"04",X"02",X"00",
    X"00",X"00",X"63",X"00",X"41",X"43",X"03",X"00",
    X"00",X"43",X"80",X"00",X"00",X"00",X"64",X"00",
    X"41",X"43",X"10",X"07",X"00",X"19",X"00",X"07",
    X"80",X"00",X"00",X"00",X"65",X"00",X"41",X"43",
    X"02",X"00",X"00",X"42",X"00",X"00",X"00",X"66",
    X"00",X"41",X"43",X"10",X"06",X"00",X"19",X"00",
    X"06",X"00",X"00",X"00",X"44",X"00",X"6F",X"00",
    X"6E",X"00",X"65",X"00",X"00",X"00",X"C6",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );

begin

    uut: entity work.mips_cpu
    port map (
        interrupt   => interrupt,
        
        data_rd_addr=> rd_addr,
        data_rd_vma => vma_data,
        data_rd     => data_r,
        
        code_rd_addr=> code_addr,
        code_rd     => code_r,
        code_rd_vma => vma_code,
        
        data_wr_addr=> wr_addr,
        data_wr     => data_w,
        byte_we     => byte_we,

        mem_wait    => mem_wait,
        
        clk         => clk,
        reset       => reset
    );

    ---------------------------------------------------------------------------
    -- Master clock: free running clock used as main module clock
    run_master_clock:
    process(done, clk)
    begin
        if done = '0' then
            clk <= not clk after T/2;
        end if;
    end process run_master_clock;

    drive_uut:
    process
    variable l : line;
    begin
        wait for T*4;
        reset <= '0';
        
        wait for T*SIMULATION_LENGTH;

        -- Flush console output to log console file (in case the end of the
        -- simulation caugh an unterminated line in the buffer)
        if con_line_ix > 1 then
            write(l, con_line_buf(1 to con_line_ix));
            writeline(con_file, l);
        end if;

        print("TB0 finished");
        done <= '1';
        wait;
        
    end process drive_uut;
    
    mem_wait <= '0'; -- memory wait input not simulated in this test bench
    

    -- RAM vs. IO data read mux
    data_r <= data_ram when prev_rd_addr(31 downto 28)/=X"2" else data_uart;
    
    -- UART read registers; only status, and hardwired, for the time being
    data_uart <= data_uart_status;
    data_uart_status <= X"0000000" & "00" & uart_tx_rdy & uart_rx_rdy;


    -- 'full' read address, used for simulation display only
    full_rd_addr <= rd_addr;
    full_wr_addr <= wr_addr & "00";
    full_code_addr <= code_addr & "00";

    data_addr_rd <= full_rd_addr(ADDR_SIZE-1+2 downto 2);
    addr_wr <= full_wr_addr(ADDR_SIZE-1+2 downto 2);
    code_addr_rd <= full_code_addr(ADDR_SIZE-1+2 downto 2);


    write_process:
    process(clk)
    variable i : integer;
    variable uart_data : integer;
    begin
        if clk'event and clk='1' then
            if reset='1' then
                data_ram <= (others =>'0');
            else
                prev_rd_addr <= rd_addr;
                
                data_ram <= 
                  ram3(conv_integer(unsigned(data_addr_rd))) &
                  ram2(conv_integer(unsigned(data_addr_rd))) &
                  ram1(conv_integer(unsigned(data_addr_rd))) &
                  ram0(conv_integer(unsigned(data_addr_rd)));
                  
                code_r <= 
                  ram3(conv_integer(unsigned(code_addr_rd))) &
                  ram2(conv_integer(unsigned(code_addr_rd))) &
                  ram1(conv_integer(unsigned(code_addr_rd))) &
                  ram0(conv_integer(unsigned(code_addr_rd)));
            end if;
            
            if byte_we/="0000" then
                if full_wr_addr(31 downto 28)=X"2" then
                    -- Write to UART
                    
                    -- If we're simulating the UART TX time, pulse RDY low
                    if SIMULATED_UART_TX_TIME > 0 us then
                        uart_tx_rdy <= '0', '1' after SIMULATED_UART_TX_TIME;
                    end if;
                    
                    -- TX data may come from the high or low byte (opcodes.s
                    -- uses high byte, no_op.c uses low)
                    if byte_we(0)='1' then
                        uart_data := conv_integer(unsigned(data_w(7 downto 0)));
                    else
                        uart_data := conv_integer(unsigned(data_w(31 downto 24)));
                    end if;
                    
                    -- UART TX data goes to output after a bit of line-buffering
                    -- and editing
                    if uart_data = 10 then
                        -- CR received: print output string and clear it
                        print(con_file, con_line_buf(1 to con_line_ix));
                        con_line_ix <= 1;
                        for i in 1 to con_line_buf'high loop
                           con_line_buf(i) <= ' ';
                        end loop;
                    elsif uart_data = 13 then
                        -- ignore LF
                    else
                        -- append char to output string
                        if con_line_ix < con_line_buf'high then
                            con_line_buf(con_line_ix) <= character'val(uart_data);
                            con_line_ix <= con_line_ix + 1;
                        end if;
                    end if;
                else
                    -- Write to RAM
                    if byte_we(3)='1' then
                        ram3(conv_integer(unsigned(addr_wr))) <= data_w(31 downto 24);
                    end if;
                    if byte_we(2)='1' then
                        ram2(conv_integer(unsigned(addr_wr))) <= data_w(23 downto 16);
                    end if;
                    if byte_we(1)='1' then
                        ram1(conv_integer(unsigned(addr_wr))) <= data_w(15 downto  8);
                    end if;
                    if byte_we(0)='1' then
                        ram0(conv_integer(unsigned(addr_wr))) <= data_w( 7 downto  0);
                    end if;
                end if;
            end if;
        end if;
    end process write_process;
                  
    log_execution:
    process
    begin
        log_cpu_activity(clk, reset, done, 
                         "mips_tb1/uut", log_info, "log_info", log_file);
        wait;
    end process log_execution;
                  
                  
--    signalspy_rbank:
--    process
--    begin
--        init_signal_spy("/mips_tb1/uut/p1_rbank", "rbank", 0, -1);
--        init_signal_spy("/mips_tb1/uut/p0_pc_reg", "pc", 0, -1);
--        init_signal_spy("/mips_tb1/uut/mult_div/upper_reg", "reg_hi", 0, -1);
--        init_signal_spy("/mips_tb1/uut/mult_div/lower_reg", "reg_lo", 0, -1);
--        init_signal_spy("/mips_tb1/uut/mult_div/negate_reg", "negate_reg_lo", 0, -1);
--        init_signal_spy("/mips_tb1/uut/cp0_epc", "cp0_epc", 0, -1);
--        init_signal_spy("/mips_tb1/uut/p2_ld_upper_byte", "ld_upper_byte", 0, -1);
--        init_signal_spy("/mips_tb1/uut/p2_ld_upper_byte", "ld_upper_hword", 0, -1);
--        wait;
--    end process signalspy_rbank;
--
--    log_cpu_activity:
--    process(clk)
--    variable prev_rbank : t_rbank := (others => X"00000000");
--    variable ri : std_logic_vector(7 downto 0);
--    variable full_pc : t_word := (others => '0');
--    variable prev_pc : t_word := (others => '0');
--    variable prev_hi : t_word := (others => '0');
--    variable prev_lo : t_word := (others => '0');
--    variable prev_epc : std_logic_vector(31 downto 2) := (others => '0');
--    variable wr_data : t_word := (others => '0');
--    variable temp : t_word := (others => '0');
--    variable size : std_logic_vector(7 downto 0) := X"00";
--    variable prev_vma_data : std_logic := '0';
--    variable prev_rd_addr : t_word := (others => '0');
--    variable rd_size : std_logic_vector(7 downto 0) := X"00";
--    begin
--        -- we'll be sampling control & data signals at falling edge, when 
--        -- they're stable
--        if clk'event and clk='0' then
--            if reset='0' then
--            
--                -- log memory loads (data only)
--                -- IMPORTANT: memory reads should be logged first because we're
--                -- logging them the cycle after they actually happen. If you put
--                -- the log code after any other log, the order of the operations 
--                -- will appear wrong in the log even though it is not.
--                if prev_vma_data='1' then
--                    if ld_upper_hword='1' then
--                        rd_size := X"04";
--                    elsif ld_upper_byte='1' then
--                        rd_size := X"02";
--                    else
--                        rd_size := X"01";
--                    end if;
--                    print(l_file, "("& hstr(prev_pc) &") ["& hstr(prev_rd_addr) &"] <"&
--                          "**"&
--                          --hstr(rd_size)& 
--                          ">="& hstr(data_r)& " RD");
--                end if;
--                prev_vma_data := vma_data;
--                prev_rd_addr := full_rd_addr;
--                
--                -- log register changes
--                ri := X"00";
--                for i in 0 to 31 loop
--                    if prev_rbank(i)/=rbank(i) then
--                        print(l_file, "("& hstr(full_pc)& ") ["& hstr(ri)& "]="& hstr(rbank(i)));
--                    end if;
--                    ri := ri + 1;
--                end loop;
--
--                -- log aux register changes, only when pipeline is not stalled
--                if prev_lo /= reg_lo and reg_lo(0)/='U' and vma_code='1' then
--                    -- we're observing the value of reg_lo, but the mult core
--                    -- will output the negated value in some cases. We
--                    -- have to mimic that behavior.
--                    if negate_reg_lo='1' then
--                        -- negate reg_lo before displaying
--                        prev_lo := not reg_lo;
--                        prev_lo := prev_lo + 1;
--                        print(l_file, "("& hstr(full_pc)& ") [LO]="& hstr(prev_lo));
--                    else
--                        print(l_file, "("& hstr(full_pc)& ") [LO]="& hstr(reg_lo));
--                    end if;
--                end if;
--                if prev_hi /= reg_hi and reg_hi(0)/='U' and vma_code='1' then
--                    print(l_file, "("& hstr(full_pc)& ") [HI]="& hstr(reg_hi));
--                end if;                
--                if prev_epc /= cp0_epc and cp0_epc(31)/='U'  then
--                    temp := cp0_epc & "00";
--                    print(l_file, "("& hstr(full_pc)& ") [EP]="& hstr(temp));
--                end if;
--
--                -- 'remember' last value of hi and lo only when pipeline is not
--                -- stalled; that's because we don't want to be tracking the
--                -- changing values when mul/div is running (because the SW 
--                -- simulator doesn't)
--                if vma_code='1' then
--                    prev_hi := reg_hi;
--                    prev_lo := reg_lo;
--                end if;
--
--
--                full_pc := pc & "00";
--                prev_pc := full_pc;
--                prev_rbank := rbank;
--                prev_epc := cp0_epc;
--                
--                -- log memory writes
--                if byte_we/="0000" then
--                    wr_data := X"00000000";
--                    if byte_we(3)='1' then
--                        wr_data(31 downto 24) := data_w(31 downto 24);
--                    end if;
--                    if byte_we(2)='1' then
--                        wr_data(23 downto 16) := data_w(23 downto 16);
--                    end if;
--                    if byte_we(1)='1' then
--                        wr_data(15 downto  8) := data_w(15 downto  8);
--                    end if;
--                    if byte_we(0)='1' then
--                        wr_data( 7 downto  0) := data_w( 7 downto  0);
--                    end if;
--                    size := "0000" & byte_we; -- mask, really
--                    print(l_file, "("& hstr(full_pc) &") ["& hstr(full_wr_addr) &"] |"& hstr(size)& "|="& hstr(wr_data)& " WR" );
--                end if;
--
--            end if;
--        end if;
--    end process log_cpu_activity;

end testbench;
