--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- This file contains object code in the form of a VHDL byte table constant.
-- This constant can be used to initialize FPGA memories for synthesis or
-- simulation.
-- Note that the object code is stored as a plain byte table in byte address
-- order. This table knows nothing of data endianess and can be used to
-- initialize 32-, 16- or 8-bit-wide memory -- memory initialization functions
-- can be found in package mips_pkg.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mips_pkg.all;

package obj_code_pkg is

constant obj_code : t_obj_code(0 to 3678) := (
  X"10", X"00", X"00", X"7c", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"40", X"1a", X"68", X"00", X"00", X"1a", X"d0", X"82", 
  X"33", X"5a", X"00", X"1f", X"34", X"1b", X"00", X"08", 
  X"13", X"5b", X"00", X"09", X"23", X"7b", X"00", X"01", 
  X"13", X"5b", X"00", X"05", X"23", X"7b", X"00", X"01", 
  X"17", X"5b", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"a2", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"40", X"1b", X"70", X"00", X"40", X"1a", X"68", X"00", 
  X"00", X"1a", X"d7", X"c2", X"33", X"5a", X"00", X"01", 
  X"17", X"40", X"00", X"03", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"42", X"00", X"00", X"10", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"fe", X"40", X"84", X"60", X"00", 
  X"0f", X"f0", X"00", X"86", X"00", X"00", X"00", X"00", 
  X"3c", X"04", X"bf", X"c0", X"24", X"84", X"06", X"b4", 
  X"00", X"80", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"3c", X"05", X"00", X"01", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"ff", X"00", X"85", X"28", X"25", 
  X"40", X"85", X"60", X"00", X"24", X"04", X"00", X"00", 
  X"24", X"06", X"00", X"00", X"24", X"05", X"00", X"ff", 
  X"ac", X"86", X"00", X"00", X"00", X"c5", X"08", X"2a", 
  X"14", X"20", X"ff", X"fd", X"20", X"c6", X"00", X"01", 
  X"24", X"04", X"00", X"00", X"24", X"06", X"00", X"00", 
  X"24", X"05", X"00", X"ff", X"8c", X"80", X"00", X"00", 
  X"20", X"84", X"00", X"10", X"00", X"c5", X"08", X"2a", 
  X"14", X"20", X"ff", X"fc", X"20", X"c6", X"00", X"01", 
  X"3c", X"05", X"00", X"02", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"ff", X"00", X"85", X"28", X"25", 
  X"03", X"e0", X"00", X"08", X"40", X"85", X"60", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"3c", X"1b", X"00", X"00", X"27", X"7b", X"00", X"3c", 
  X"af", X"7d", X"ff", X"f0", X"af", X"7f", X"ff", X"ec", 
  X"af", X"68", X"ff", X"e8", X"af", X"69", X"ff", X"e4", 
  X"af", X"6a", X"ff", X"e0", X"03", X"60", X"e8", X"21", 
  X"40", X"08", X"70", X"00", X"8d", X"1a", X"00", X"00", 
  X"40", X"1b", X"68", X"00", X"07", X"70", X"00", X"2d", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"4e", X"82", 
  X"39", X"28", X"00", X"1f", X"11", X"00", X"00", X"1f", 
  X"39", X"28", X"00", X"1c", X"11", X"00", X"00", X"13", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"8f", X"aa", X"ff", X"e0", 
  X"8f", X"a9", X"ff", X"e4", X"8f", X"a8", X"ff", X"e8", 
  X"8f", X"bf", X"ff", X"ec", X"8f", X"bd", X"ff", X"f0", 
  X"40", X"1b", X"70", X"00", X"40", X"1a", X"68", X"00", 
  X"00", X"1a", X"d7", X"c2", X"33", X"5a", X"00", X"01", 
  X"17", X"40", X"00", X"03", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"42", X"00", X"00", X"10", X"33", X"5b", X"00", X"3f", 
  X"3b", X"68", X"00", X"20", X"11", X"00", X"00", X"14", 
  X"3b", X"68", X"00", X"21", X"11", X"00", X"00", X"1c", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"0b", X"f0", X"00", X"b7", 
  X"00", X"00", X"00", X"00", X"33", X"5b", X"00", X"3f", 
  X"3b", X"68", X"00", X"00", X"11", X"00", X"00", X"1e", 
  X"3b", X"68", X"00", X"04", X"11", X"00", X"00", X"29", 
  X"00", X"00", X"00", X"00", X"3c", X"08", X"20", X"01", 
  X"ad", X"1a", X"04", X"00", X"0b", X"f0", X"00", X"b7", 
  X"00", X"00", X"00", X"00", X"8d", X"1a", X"00", X"04", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"0f", X"f0", X"01", X"61", X"3c", X"0a", X"80", X"00", 
  X"00", X"00", X"40", X"21", X"03", X"6a", X"48", X"24", 
  X"15", X"20", X"00", X"03", X"00", X"0a", X"50", X"42", 
  X"15", X"40", X"ff", X"fc", X"25", X"08", X"00", X"01", 
  X"0b", X"f0", X"01", X"17", X"01", X"00", X"d8", X"21", 
  X"0f", X"f0", X"01", X"61", X"3c", X"0a", X"80", X"00", 
  X"00", X"00", X"40", X"21", X"03", X"6a", X"48", X"24", 
  X"11", X"20", X"00", X"03", X"00", X"0a", X"50", X"42", 
  X"15", X"40", X"ff", X"fc", X"25", X"08", X"00", X"01", 
  X"0b", X"f0", X"01", X"17", X"01", X"00", X"d8", X"21", 
  X"0f", X"f0", X"01", X"61", X"00", X"00", X"00", X"00", 
  X"00", X"1a", X"41", X"82", X"31", X"08", X"00", X"1f", 
  X"00", X"1a", X"4a", X"c2", X"31", X"29", X"00", X"1f", 
  X"01", X"09", X"50", X"21", X"00", X"0a", X"50", X"23", 
  X"25", X"4a", X"00", X"1f", X"01", X"5b", X"d8", X"04", 
  X"01", X"5b", X"d8", X"06", X"0b", X"f0", X"01", X"17", 
  X"01", X"1b", X"d8", X"06", X"0f", X"f0", X"01", X"61", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"41", X"82", 
  X"31", X"08", X"00", X"1f", X"00", X"1a", X"4a", X"c2", 
  X"31", X"29", X"00", X"1f", X"01", X"28", X"48", X"23", 
  X"00", X"09", X"58", X"23", X"25", X"6b", X"00", X"1f", 
  X"01", X"1b", X"48", X"04", X"3c", X"0a", X"ff", X"ff", 
  X"35", X"4a", X"ff", X"ff", X"01", X"6a", X"50", X"04", 
  X"01", X"6a", X"50", X"06", X"01", X"0a", X"50", X"04", 
  X"01", X"2a", X"48", X"24", X"01", X"40", X"50", X"27", 
  X"0f", X"f0", X"01", X"61", X"00", X"1a", X"d1", X"40", 
  X"00", X"1a", X"d1", X"42", X"03", X"6a", X"d8", X"24", 
  X"03", X"69", X"d8", X"25", X"0b", X"f0", X"01", X"17", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"4c", X"02", 
  X"31", X"29", X"00", X"1f", X"3c", X"08", X"bf", X"c0", 
  X"25", X"08", X"04", X"84", X"00", X"09", X"48", X"c0", 
  X"01", X"09", X"40", X"20", X"01", X"00", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"00", X"b7", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"60", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"61", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"62", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"63", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"64", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"65", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"66", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"67", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"af", X"bb", X"ff", X"e8", X"0b", X"f0", X"01", X"1f", 
  X"af", X"bb", X"ff", X"e4", X"0b", X"f0", X"01", X"1f", 
  X"af", X"bb", X"ff", X"e0", X"0b", X"f0", X"01", X"1f", 
  X"37", X"6b", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"6c", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"6d", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"6e", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"6f", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"70", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"71", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"72", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"73", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"74", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"75", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"76", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"77", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"78", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"79", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"7a", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"7b", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"37", X"7c", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"af", X"bb", X"ff", X"ec", X"0b", X"f0", X"01", X"1f", 
  X"37", X"7e", X"00", X"00", X"0b", X"f0", X"01", X"1f", 
  X"af", X"bb", X"ff", X"f0", X"af", X"bf", X"00", X"00", 
  X"00", X"1a", X"dd", X"42", X"33", X"7b", X"00", X"1f", 
  X"3c", X"08", X"bf", X"c0", X"25", X"08", X"05", X"b4", 
  X"00", X"1b", X"d8", X"c0", X"01", X"1b", X"40", X"20", 
  X"01", X"00", X"f8", X"09", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"34", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e8", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e4", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"e0", X"03", X"e0", X"00", X"08", 
  X"35", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"35", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"9b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"bb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"36", X"fb", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"1b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"3b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"5b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"7b", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"37", X"9a", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"f0", X"03", X"e0", X"00", X"08", 
  X"37", X"db", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"8f", X"bb", X"ff", X"ec", X"3c", X"1c", X"00", X"00", 
  X"27", X"9c", X"7f", X"f0", X"3c", X"05", X"00", X"00", 
  X"24", X"a5", X"00", X"00", X"3c", X"04", X"00", X"00", 
  X"24", X"84", X"00", X"00", X"3c", X"1d", X"00", X"00", 
  X"27", X"bd", X"04", X"28", X"ac", X"a0", X"00", X"00", 
  X"00", X"a4", X"18", X"2a", X"14", X"60", X"ff", X"fd", 
  X"24", X"a5", X"00", X"04", X"3c", X"04", X"00", X"00", 
  X"24", X"84", X"00", X"00", X"3c", X"05", X"bf", X"c0", 
  X"24", X"a5", X"0e", X"60", X"10", X"a4", X"00", X"0b", 
  X"00", X"00", X"00", X"00", X"3c", X"10", X"00", X"00", 
  X"26", X"10", X"00", X"00", X"12", X"00", X"00", X"07", 
  X"00", X"00", X"00", X"00", X"8c", X"a8", X"00", X"00", 
  X"24", X"a5", X"00", X"04", X"ac", X"88", X"00", X"00", 
  X"24", X"84", X"00", X"04", X"16", X"00", X"ff", X"fb", 
  X"26", X"10", X"ff", X"fc", X"0f", X"f0", X"01", X"cd", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"01", X"cb", 
  X"00", X"00", X"00", X"00", X"3c", X"04", X"bf", X"c0", 
  X"27", X"bd", X"ff", X"e8", X"af", X"bf", X"00", X"14", 
  X"0f", X"f0", X"03", X"40", X"24", X"84", X"0e", X"04", 
  X"3c", X"04", X"bf", X"c0", X"0f", X"f0", X"03", X"40", 
  X"24", X"84", X"0e", X"2c", X"3c", X"04", X"bf", X"c0", 
  X"8f", X"bf", X"00", X"14", X"24", X"84", X"0e", X"44", 
  X"0b", X"f0", X"03", X"40", X"27", X"bd", X"00", X"18", 
  X"10", X"80", X"00", X"09", X"00", X"00", X"00", X"00", 
  X"8c", X"82", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"a0", X"45", X"00", X"00", X"8c", X"82", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"24", X"42", X"00", X"01", 
  X"03", X"e0", X"00", X"08", X"ac", X"82", X"00", X"00", 
  X"0b", X"f0", X"03", X"6e", X"00", X"a0", X"20", X"21", 
  X"27", X"bd", X"ff", X"d8", X"af", X"b2", X"00", X"18", 
  X"af", X"b1", X"00", X"14", X"af", X"b0", X"00", X"10", 
  X"af", X"bf", X"00", X"24", X"af", X"b4", X"00", X"20", 
  X"af", X"b3", X"00", X"1c", X"00", X"c0", X"90", X"21", 
  X"00", X"80", X"88", X"21", X"18", X"c0", X"00", X"32", 
  X"00", X"a0", X"80", X"21", X"90", X"a2", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"00", X"3d", 
  X"00", X"a0", X"10", X"21", X"00", X"00", X"18", X"21", 
  X"24", X"42", X"00", X"01", X"90", X"44", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"14", X"80", X"ff", X"fc", 
  X"24", X"63", X"00", X"01", X"00", X"72", X"10", X"2a", 
  X"14", X"40", X"00", X"02", X"02", X"43", X"90", X"23", 
  X"00", X"00", X"90", X"21", X"30", X"e2", X"00", X"02", 
  X"10", X"40", X"00", X"22", X"30", X"e7", X"00", X"01", 
  X"10", X"e0", X"00", X"22", X"24", X"14", X"00", X"30", 
  X"00", X"00", X"98", X"21", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"a0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"02", X"20", X"20", X"21", 
  X"0f", X"f0", X"01", X"da", X"26", X"10", X"00", X"01", 
  X"92", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"14", X"a0", X"ff", X"fa", X"26", X"73", X"00", X"01", 
  X"1a", X"40", X"00", X"08", X"02", X"40", X"80", X"21", 
  X"26", X"10", X"ff", X"ff", X"02", X"20", X"20", X"21", 
  X"0f", X"f0", X"01", X"da", X"02", X"80", X"28", X"21", 
  X"16", X"00", X"ff", X"fc", X"26", X"10", X"ff", X"ff", 
  X"02", X"72", X"98", X"21", X"8f", X"bf", X"00", X"24", 
  X"02", X"60", X"10", X"21", X"8f", X"b4", X"00", X"20", 
  X"8f", X"b3", X"00", X"1c", X"8f", X"b2", X"00", X"18", 
  X"8f", X"b1", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"30", X"e7", X"00", X"01", X"14", X"e0", X"ff", X"e0", 
  X"24", X"14", X"00", X"20", X"1a", X"40", X"ff", X"de", 
  X"02", X"40", X"98", X"21", X"26", X"73", X"ff", X"ff", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"01", X"da", 
  X"02", X"80", X"28", X"21", X"16", X"60", X"ff", X"fc", 
  X"26", X"73", X"ff", X"ff", X"26", X"73", X"00", X"01", 
  X"02", X"40", X"98", X"21", X"0b", X"f0", X"02", X"05", 
  X"00", X"00", X"90", X"21", X"00", X"00", X"18", X"21", 
  X"0b", X"f0", X"01", X"ff", X"02", X"43", X"90", X"23", 
  X"27", X"bd", X"ff", X"c8", X"af", X"b4", X"00", X"30", 
  X"af", X"b2", X"00", X"28", X"af", X"b1", X"00", X"24", 
  X"af", X"bf", X"00", X"34", X"af", X"b3", X"00", X"2c", 
  X"af", X"b0", X"00", X"20", X"00", X"a0", X"10", X"21", 
  X"8f", X"b4", X"00", X"48", X"8f", X"b2", X"00", X"4c", 
  X"10", X"a0", X"00", X"3f", X"00", X"80", X"88", X"21", 
  X"14", X"e0", X"00", X"31", X"24", X"03", X"00", X"0a", 
  X"00", X"00", X"38", X"21", X"10", X"40", X"00", X"49", 
  X"a3", X"a0", X"00", X"1b", X"8f", X"a5", X"00", X"50", 
  X"27", X"b3", X"00", X"1b", X"24", X"a5", X"ff", X"c6", 
  X"14", X"c0", X"00", X"02", X"00", X"46", X"00", X"1b", 
  X"00", X"07", X"00", X"0d", X"00", X"00", X"18", X"10", 
  X"28", X"64", X"00", X"0a", X"00", X"00", X"00", X"00", 
  X"14", X"c0", X"00", X"02", X"00", X"46", X"00", X"1b", 
  X"00", X"07", X"00", X"0d", X"00", X"00", X"10", X"12", 
  X"14", X"80", X"00", X"02", X"26", X"73", X"ff", X"ff", 
  X"00", X"65", X"18", X"21", X"24", X"63", X"00", X"30", 
  X"14", X"40", X"ff", X"f1", X"a2", X"63", X"00", X"00", 
  X"14", X"e0", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"80", X"21", X"02", X"20", X"20", X"21", 
  X"02", X"60", X"28", X"21", X"02", X"80", X"30", X"21", 
  X"0f", X"f0", X"01", X"e6", X"02", X"40", X"38", X"21", 
  X"8f", X"bf", X"00", X"34", X"00", X"50", X"10", X"21", 
  X"8f", X"b4", X"00", X"30", X"8f", X"b3", X"00", X"2c", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"12", X"80", X"00", X"0f", 
  X"32", X"42", X"00", X"02", X"10", X"40", X"00", X"0d", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"01", X"da", 
  X"24", X"05", X"00", X"2d", X"26", X"94", X"ff", X"ff", 
  X"0b", X"f0", X"02", X"5b", X"24", X"10", X"00", X"01", 
  X"14", X"c3", X"ff", X"d0", X"00", X"00", X"38", X"21", 
  X"04", X"a1", X"ff", X"ce", X"00", X"00", X"00", X"00", 
  X"00", X"05", X"10", X"23", X"0b", X"f0", X"02", X"43", 
  X"24", X"07", X"00", X"01", X"26", X"73", X"ff", X"ff", 
  X"24", X"02", X"00", X"2d", X"a2", X"62", X"00", X"00", 
  X"0b", X"f0", X"02", X"5b", X"00", X"00", X"80", X"21", 
  X"27", X"a5", X"00", X"10", X"02", X"80", X"30", X"21", 
  X"02", X"40", X"38", X"21", X"24", X"02", X"00", X"30", 
  X"a3", X"a2", X"00", X"10", X"0f", X"f0", X"01", X"e6", 
  X"a3", X"a0", X"00", X"11", X"8f", X"bf", X"00", X"34", 
  X"8f", X"b4", X"00", X"30", X"8f", X"b3", X"00", X"2c", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"10", X"e0", X"ff", X"cc", 
  X"27", X"b3", X"00", X"1b", X"0b", X"f0", X"02", X"69", 
  X"00", X"00", X"00", X"00", X"27", X"bd", X"ff", X"b8", 
  X"af", X"b4", X"00", X"38", X"af", X"b0", X"00", X"28", 
  X"af", X"bf", X"00", X"44", X"af", X"b6", X"00", X"40", 
  X"af", X"b5", X"00", X"3c", X"af", X"b3", X"00", X"34", 
  X"af", X"b2", X"00", X"30", X"af", X"b1", X"00", X"2c", 
  X"00", X"a0", X"80", X"21", X"90", X"a5", X"00", X"00", 
  X"00", X"80", X"a0", X"21", X"10", X"a0", X"00", X"a0", 
  X"af", X"a6", X"00", X"50", X"00", X"00", X"90", X"21", 
  X"24", X"13", X"00", X"25", X"24", X"15", X"00", X"2d", 
  X"24", X"11", X"00", X"30", X"3c", X"16", X"bf", X"c0", 
  X"14", X"b3", X"00", X"53", X"00", X"00", X"00", X"00", 
  X"26", X"10", X"00", X"01", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"a0", X"00", X"3e", 
  X"00", X"00", X"00", X"00", X"10", X"b3", X"00", X"4c", 
  X"00", X"00", X"00", X"00", X"10", X"b5", X"00", X"54", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"18", X"21", 
  X"14", X"b1", X"00", X"07", X"24", X"a2", X"ff", X"d0", 
  X"26", X"10", X"00", X"01", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"b1", X"ff", X"fc", 
  X"34", X"63", X"00", X"02", X"24", X"a2", X"ff", X"d0", 
  X"30", X"42", X"00", X"ff", X"2c", X"42", X"00", X"0a", 
  X"10", X"40", X"00", X"0d", X"00", X"00", X"10", X"21", 
  X"00", X"02", X"20", X"40", X"00", X"02", X"10", X"c0", 
  X"00", X"82", X"10", X"21", X"26", X"10", X"00", X"01", 
  X"00", X"45", X"10", X"21", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"24", X"a4", X"ff", X"d0", 
  X"30", X"84", X"00", X"ff", X"2c", X"84", X"00", X"0a", 
  X"14", X"80", X"ff", X"f5", X"24", X"42", X"ff", X"d0", 
  X"24", X"04", X"00", X"73", X"10", X"a4", X"00", X"3c", 
  X"24", X"04", X"00", X"64", X"10", X"a4", X"00", X"46", 
  X"02", X"80", X"20", X"21", X"24", X"04", X"00", X"78", 
  X"10", X"a4", X"00", X"51", X"02", X"80", X"20", X"21", 
  X"24", X"04", X"00", X"58", X"10", X"a4", X"00", X"55", 
  X"02", X"80", X"20", X"21", X"24", X"04", X"00", X"75", 
  X"10", X"a4", X"00", X"60", X"02", X"80", X"20", X"21", 
  X"24", X"04", X"00", X"63", X"14", X"a4", X"00", X"24", 
  X"26", X"10", X"00", X"01", X"8f", X"a9", X"00", X"50", 
  X"27", X"a5", X"00", X"20", X"8d", X"28", X"00", X"00", 
  X"02", X"80", X"20", X"21", X"25", X"29", X"00", X"04", 
  X"00", X"40", X"30", X"21", X"00", X"60", X"38", X"21", 
  X"af", X"a9", X"00", X"50", X"a3", X"a8", X"00", X"20", 
  X"0f", X"f0", X"01", X"e6", X"a3", X"a0", X"00", X"21", 
  X"92", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"14", X"a0", X"ff", X"bd", X"02", X"42", X"90", X"21", 
  X"12", X"80", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"8e", X"82", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"a0", X"40", X"00", X"00", X"8f", X"bf", X"00", X"44", 
  X"02", X"40", X"10", X"21", X"8f", X"b6", X"00", X"40", 
  X"8f", X"b5", X"00", X"3c", X"8f", X"b4", X"00", X"38", 
  X"8f", X"b3", X"00", X"34", X"8f", X"b2", X"00", X"30", 
  X"8f", X"b1", X"00", X"2c", X"8f", X"b0", X"00", X"28", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"48", 
  X"0f", X"f0", X"01", X"da", X"02", X"80", X"20", X"21", 
  X"26", X"52", X"00", X"01", X"26", X"10", X"00", X"01", 
  X"92", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"14", X"a0", X"ff", X"a5", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"02", X"e8", X"00", X"00", X"00", X"00", 
  X"26", X"10", X"00", X"01", X"92", X"05", X"00", X"00", 
  X"0b", X"f0", X"02", X"b0", X"24", X"03", X"00", X"01", 
  X"8f", X"a4", X"00", X"50", X"00", X"00", X"00", X"00", 
  X"8c", X"85", X"00", X"00", X"24", X"84", X"00", X"04", 
  X"10", X"a0", X"00", X"31", X"af", X"a4", X"00", X"50", 
  X"02", X"80", X"20", X"21", X"00", X"40", X"30", X"21", 
  X"0f", X"f0", X"01", X"e6", X"00", X"60", X"38", X"21", 
  X"0b", X"f0", X"02", X"fb", X"02", X"42", X"90", X"21", 
  X"8f", X"a8", X"00", X"50", X"00", X"00", X"00", X"00", 
  X"8d", X"05", X"00", X"00", X"24", X"06", X"00", X"0a", 
  X"25", X"08", X"00", X"04", X"24", X"07", X"00", X"01", 
  X"af", X"a2", X"00", X"10", X"24", X"02", X"00", X"61", 
  X"af", X"a8", X"00", X"50", X"af", X"a3", X"00", X"14", 
  X"0f", X"f0", X"02", X"34", X"af", X"a2", X"00", X"18", 
  X"0b", X"f0", X"02", X"fb", X"02", X"42", X"90", X"21", 
  X"8f", X"a8", X"00", X"50", X"00", X"00", X"00", X"00", 
  X"8d", X"05", X"00", X"00", X"24", X"06", X"00", X"10", 
  X"25", X"08", X"00", X"04", X"0b", X"f0", X"03", X"18", 
  X"00", X"00", X"38", X"21", X"8f", X"a8", X"00", X"50", 
  X"00", X"00", X"00", X"00", X"8d", X"05", X"00", X"00", 
  X"24", X"06", X"00", X"10", X"25", X"08", X"00", X"04", 
  X"af", X"a2", X"00", X"10", X"00", X"00", X"38", X"21", 
  X"24", X"02", X"00", X"41", X"af", X"a8", X"00", X"50", 
  X"af", X"a3", X"00", X"14", X"0f", X"f0", X"02", X"34", 
  X"af", X"a2", X"00", X"18", X"0b", X"f0", X"02", X"fb", 
  X"02", X"42", X"90", X"21", X"8f", X"a8", X"00", X"50", 
  X"00", X"00", X"00", X"00", X"8d", X"05", X"00", X"00", 
  X"24", X"06", X"00", X"0a", X"25", X"08", X"00", X"04", 
  X"0b", X"f0", X"03", X"18", X"00", X"00", X"38", X"21", 
  X"0b", X"f0", X"03", X"0c", X"26", X"c5", X"0e", X"58", 
  X"0b", X"f0", X"02", X"e8", X"00", X"00", X"90", X"21", 
  X"27", X"bd", X"ff", X"e0", X"27", X"a2", X"00", X"24", 
  X"00", X"80", X"18", X"21", X"af", X"a5", X"00", X"24", 
  X"af", X"a6", X"00", X"28", X"00", X"00", X"20", X"21", 
  X"00", X"60", X"28", X"21", X"00", X"40", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"af", X"a7", X"00", X"2c", 
  X"0f", X"f0", X"02", X"91", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"27", X"a2", X"00", X"28", 
  X"af", X"a4", X"00", X"20", X"af", X"a6", X"00", X"28", 
  X"27", X"a4", X"00", X"20", X"00", X"40", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"af", X"a7", X"00", X"2c", 
  X"0f", X"f0", X"02", X"91", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"27", X"a2", X"00", X"2c", 
  X"af", X"a4", X"00", X"20", X"00", X"c0", X"28", X"21", 
  X"27", X"a4", X"00", X"20", X"00", X"40", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"af", X"a7", X"00", X"2c", 
  X"0f", X"f0", X"02", X"91", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"00", X"80", X"10", X"21", X"3c", X"05", X"20", X"00", 
  X"8c", X"a3", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"30", X"63", X"00", X"02", X"10", X"60", X"ff", X"fc", 
  X"3c", X"03", X"20", X"00", X"ac", X"62", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"3c", X"03", X"20", X"00", X"8c", X"62", X"00", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"42", X"00", X"01", 
  X"10", X"40", X"ff", X"fc", X"3c", X"02", X"20", X"00", 
  X"8c", X"42", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"02", X"16", X"02", X"63", X"6f", X"6d", X"70", 
  X"69", X"6c", X"65", X"20", X"74", X"69", X"6d", X"65", 
  X"3a", X"20", X"4a", X"75", X"6e", X"20", X"20", X"39", 
  X"20", X"32", X"30", X"31", X"32", X"20", X"2d", X"2d", 
  X"20", X"31", X"36", X"3a", X"33", X"38", X"3a", X"30", 
  X"32", X"0a", X"00", X"00", X"67", X"63", X"63", X"20", 
  X"76", X"65", X"72", X"73", X"69", X"6f", X"6e", X"3a", 
  X"20", X"20", X"34", X"2e", X"35", X"2e", X"32", X"0a", 
  X"00", X"00", X"00", X"00", X"0a", X"0a", X"48", X"65", 
  X"6c", X"6c", X"6f", X"20", X"57", X"6f", X"72", X"6c", 
  X"64", X"21", X"0a", X"0a", X"0a", X"00", X"00", X"00", 
  X"28", X"6e", X"75", X"6c", X"6c", X"29", X"00" 
);


end package obj_code_pkg;
