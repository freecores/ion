--##############################################################################
-- This file was generated automatically from '/src/mips_tb2_template.vhdl'.
-- 
--------------------------------------------------------------------------------
-- Simulation test bench TB2 -- not synthesizable.
--
-- Simulates the CPU core connected to a simulated external static RAM and an
-- internal BRAM block through a stub (i.e. empty).
-- BRAM is initialized with the program object code, and SRAM is initialized 
-- with data secions from program. 
-- The makefile for the source samples include targets to build simulation test 
-- benches using this template, use them as usage examples.
--
-- The memory setup is meant to test the basic 'dummy' cache. 
-- 
-- Console output (at addresses compatible to Plasma's) is logged to text file
-- "hw_sim_console_log.txt".
-- IMPORTANT: The code that echoes UART TX data to the simulation console does
-- line buffering; it will not print anything until it gets a CR (0x0d), and
-- will ifnore LFs (0x0a). Bear this in mind if you see no output when you 
-- expect it.
--
-- WARNING: Will only work on Modelsim; uses custom library SignalSpy.
--##############################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use std.textio.all;

use work.mips_pkg.all;
use work.mips_tb_pkg.all;
use work.txt_util.all;

entity mips_tb2 is
end;


architecture testbench of mips_tb2 is

-------------------------------------------------------------------------------
-- Simulation parameters

-- Master clock period
constant T : time           := 20 ns;
-- Time the UART is unavailable after writing to the TX register
-- WARNING: slite does not simulate this. The logs may be different when > 0.0!
constant SIMULATED_UART_TX_TIME : time := 0.0 us;

-- Simulation length in clock cycles, should be long enough (you have to try...)
constant SIMULATION_LENGTH : integer := 400000;

-- Simulated external SRAM size in 32-bit words 
constant SRAM_SIZE : integer := 1024;
-- Ext. SRAM address length (memory is 16 bits wide so it needs an extra address bit)
constant SRAM_ADDR_SIZE : integer := log2(SRAM_SIZE)+1;


-- BRAM table and interface signals --------------------------------------------
constant BRAM_SIZE : integer := 2048;
constant BRAM_ADDR_SIZE : integer := 11;
subtype t_bram_address is std_logic_vector(BRAM_ADDR_SIZE-1 downto 0);
-- (this table holds one byte-slice; the RAM will have 4 of these)
type t_bram is array(0 to BRAM_SIZE-1) of std_logic_vector(7 downto 0);

signal bram_rd_addr :       t_bram_address; 
signal bram_wr_addr :       t_bram_address;
signal bram_rd_data :       t_word;
signal bram_wr_data :       t_word;
signal bram_byte_we :       std_logic_vector(3 downto 0);
signal bram_data_rd_vma :   std_logic;

-- bram0 is LSB, bram3 is MSB
signal bram3 : t_bram := (
    X"10",X"00",X"40",X"0F",X"00",X"3C",X"24",X"0F",
    X"00",X"24",X"24",X"0F",X"00",X"3C",X"24",X"0F",
    X"00",X"24",X"24",X"24",X"24",X"01",X"AD",X"8D",
    X"21",X"AD",X"00",X"8D",X"00",X"21",X"AD",X"00",
    X"8D",X"00",X"8D",X"11",X"00",X"AD",X"8D",X"15",
    X"00",X"01",X"15",X"25",X"10",X"00",X"10",X"00",
    X"10",X"00",X"3C",X"24",X"0F",X"00",X"21",X"01",
    X"23",X"24",X"0F",X"00",X"3C",X"24",X"0F",X"00",
    X"24",X"20",X"AC",X"00",X"14",X"20",X"24",X"24",
    X"3C",X"24",X"8C",X"00",X"AC",X"20",X"20",X"14",
    X"20",X"3C",X"24",X"0F",X"00",X"24",X"0F",X"34",
    X"24",X"00",X"00",X"00",X"3C",X"24",X"0F",X"00",
    X"3C",X"00",X"00",X"00",X"3C",X"24",X"0F",X"00",
    X"0B",X"00",X"AF",X"23",X"3C",X"24",X"3C",X"24",
    X"00",X"00",X"8F",X"03",X"23",X"00",X"00",X"00",
    X"AF",X"23",X"01",X"24",X"0F",X"00",X"3C",X"24",
    X"0F",X"00",X"24",X"8D",X"0F",X"24",X"3C",X"24",
    X"0F",X"21",X"23",X"17",X"00",X"3C",X"24",X"0F",
    X"00",X"21",X"15",X"00",X"3C",X"24",X"0F",X"21",
    X"00",X"8F",X"03",X"23",X"3C",X"40",X"24",X"24",
    X"24",X"AC",X"00",X"14",X"20",X"40",X"3C",X"00",
    X"03",X"40",X"3C",X"80",X"10",X"24",X"8C",X"30",
    X"10",X"00",X"AC",X"10",X"00",X"03",X"00",X"3C",
    X"3C",X"24",X"20",X"00",X"00",X"00",X"30",X"00",
    X"82",X"8C",X"30",X"10",X"00",X"AC",X"14",X"20",
    X"03",X"00",X"30",X"34",X"38",X"63",X"0A",X"61",
    X"6E",X"78",X"6E",X"6D",X"72",X"74",X"00",X"6E",
    X"52",X"74",X"61",X"20",X"20",X"20",X"0A",X"20",
    X"74",X"72",X"21",X"62",X"72",X"62",X"21",X"0A",
    X"6D",X"67",X"65",X"72",X"66",X"77",X"73",X"20",
    X"53",X"74",X"64",X"73",X"00",X"65",X"6E",X"6F",
    X"65",X"75",X"6E",X"6F",X"52",X"2E",X"69",X"6F",
    X"65",X"68",X"20",X"77",X"65",X"00",X"0D",X"20",
    X"74",X"2E",X"0D",X"6D",X"66",X"72",X"66",X"77",
    X"73",X"20",X"4D",X"74",X"69",X"69",X"7A",X"6F",
    X"0D",X"00",X"64",X"20",X"70",X"0D",X"74",X"20",
    X"63",X"6F",X"72",X"38",X"74",X"61",X"20",X"6F",
    X"28",X"53",X"0D",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal bram2 : t_bram := (
    X"00",X"00",X"80",X"F0",X"00",X"04",X"84",X"F0",
    X"00",X"04",X"05",X"F0",X"00",X"04",X"84",X"F0",
    X"00",X"08",X"0A",X"0B",X"0C",X"00",X"00",X"09",
    X"2A",X"0A",X"00",X"0B",X"00",X"4A",X"0A",X"00",
    X"0B",X"00",X"09",X"A9",X"00",X"08",X"09",X"28",
    X"00",X"4B",X"40",X"08",X"00",X"00",X"00",X"00",
    X"00",X"00",X"04",X"84",X"F0",X"00",X"04",X"00",
    X"BD",X"05",X"F0",X"00",X"04",X"84",X"F0",X"00",
    X"04",X"85",X"80",X"85",X"20",X"84",X"05",X"04",
    X"07",X"E7",X"E6",X"00",X"86",X"A5",X"E7",X"A0",
    X"84",X"04",X"84",X"F0",X"00",X"04",X"F0",X"05",
    X"04",X"00",X"80",X"00",X"04",X"84",X"F0",X"00",
    X"04",X"00",X"80",X"00",X"04",X"84",X"F0",X"00",
    X"F0",X"00",X"BF",X"BD",X"04",X"84",X"05",X"A5",
    X"A0",X"00",X"BF",X"E0",X"BD",X"00",X"80",X"A0",
    X"BF",X"BD",X"E0",X"05",X"F0",X"00",X"04",X"84",
    X"F0",X"00",X"19",X"E4",X"F0",X"05",X"04",X"84",
    X"F0",X"EF",X"39",X"20",X"00",X"04",X"84",X"F0",
    X"00",X"CE",X"C0",X"00",X"04",X"84",X"F0",X"EF",
    X"00",X"BF",X"E0",X"BD",X"04",X"84",X"04",X"06",
    X"05",X"86",X"C5",X"20",X"C6",X"04",X"05",X"A5",
    X"E0",X"84",X"06",X"82",X"40",X"84",X"C3",X"63",
    X"60",X"00",X"C2",X"00",X"00",X"E0",X"00",X"06",
    X"07",X"E7",X"A5",X"A5",X"A5",X"A4",X"42",X"E2",
    X"42",X"C3",X"63",X"60",X"00",X"C2",X"A0",X"A5",
    X"E0",X"00",X"31",X"35",X"39",X"64",X"0D",X"6E",
    X"67",X"74",X"61",X"65",X"79",X"20",X"46",X"64",
    X"41",X"6F",X"74",X"20",X"20",X"30",X"0D",X"00",
    X"20",X"72",X"0A",X"61",X"65",X"61",X"0A",X"0D",
    X"70",X"20",X"20",X"73",X"65",X"6F",X"20",X"46",
    X"48",X"20",X"72",X"20",X"0A",X"73",X"67",X"64",
    X"78",X"74",X"20",X"6D",X"41",X"2E",X"66",X"75",
    X"65",X"69",X"69",X"6F",X"64",X"0A",X"45",X"6F",
    X"65",X"0A",X"00",X"70",X"20",X"73",X"65",X"6F",
    X"20",X"58",X"20",X"65",X"6E",X"61",X"61",X"6E",
    X"00",X"3C",X"20",X"64",X"3E",X"54",X"69",X"65",
    X"75",X"6E",X"6F",X"2D",X"20",X"74",X"6D",X"72",
    X"46",X"48",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal bram1 : t_bram := (
    X"00",X"00",X"60",X"00",X"00",X"BF",X"03",X"00",
    X"00",X"00",X"00",X"00",X"00",X"BF",X"03",X"00",
    X"00",X"00",X"04",X"00",X"00",X"68",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"50",X"FF",X"04",X"00",X"00",X"00",X"00",
    X"00",X"00",X"BF",X"03",X"00",X"00",X"FF",X"E8",
    X"FF",X"00",X"00",X"00",X"BF",X"03",X"00",X"00",
    X"00",X"01",X"00",X"08",X"FF",X"00",X"00",X"00",
    X"BF",X"01",X"00",X"00",X"00",X"FF",X"00",X"FF",
    X"00",X"BF",X"04",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"F8",X"00",X"BF",X"04",X"00",X"00",
    X"B0",X"00",X"F8",X"00",X"BF",X"04",X"00",X"00",
    X"00",X"00",X"00",X"FF",X"BF",X"03",X"BF",X"02",
    X"F8",X"00",X"00",X"00",X"00",X"00",X"78",X"70",
    X"00",X"FF",X"20",X"00",X"00",X"00",X"BF",X"04",
    X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"03",
    X"00",X"00",X"FF",X"FF",X"00",X"BF",X"03",X"00",
    X"00",X"FF",X"FF",X"00",X"BF",X"04",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
    X"00",X"00",X"08",X"FF",X"00",X"60",X"00",X"20",
    X"00",X"60",X"20",X"00",X"00",X"00",X"00",X"00",
    X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"20",
    X"BF",X"03",X"FF",X"28",X"28",X"10",X"00",X"90",
    X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",
    X"00",X"00",X"32",X"36",X"61",X"65",X"53",X"6E",
    X"20",X"65",X"6C",X"6D",X"20",X"30",X"6F",X"20",
    X"4D",X"70",X"20",X"20",X"20",X"78",X"00",X"68",
    X"6D",X"6F",X"0D",X"64",X"61",X"63",X"0D",X"44",
    X"69",X"74",X"66",X"74",X"77",X"72",X"6F",X"4C",
    X"20",X"61",X"65",X"30",X"0D",X"74",X"20",X"65",
    X"65",X"69",X"66",X"20",X"4D",X"20",X"20",X"20",
    X"20",X"73",X"74",X"72",X"0A",X"0D",X"6E",X"66",
    X"73",X"0D",X"44",X"20",X"66",X"74",X"77",X"72",
    X"6F",X"52",X"61",X"72",X"69",X"6C",X"74",X"3A",
    X"3A",X"65",X"6F",X"75",X"00",X"65",X"6E",X"78",
    X"74",X"20",X"6D",X"62",X"73",X"69",X"65",X"79",
    X"4C",X"29",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal bram0 : t_bram := (
    X"01",X"00",X"00",X"9C",X"00",X"C0",X"38",X"AA",
    X"00",X"00",X"08",X"B7",X"00",X"C0",X"78",X"AA",
    X"00",X"04",X"00",X"01",X"00",X"21",X"00",X"00",
    X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
    X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"08",
    X"00",X"22",X"F7",X"00",X"05",X"00",X"03",X"00",
    X"01",X"00",X"C0",X"59",X"AA",X"00",X"FC",X"21",
    X"F0",X"08",X"B7",X"00",X"C0",X"78",X"AA",X"00",
    X"00",X"40",X"00",X"2A",X"FD",X"04",X"40",X"00",
    X"C0",X"A8",X"00",X"00",X"00",X"FC",X"04",X"FA",
    X"04",X"C0",X"2A",X"AA",X"00",X"00",X"76",X"14",
    X"00",X"00",X"09",X"00",X"C0",X"73",X"AA",X"00",
    X"00",X"00",X"09",X"00",X"C0",X"15",X"AA",X"00",
    X"68",X"00",X"00",X"FC",X"C0",X"D1",X"C0",X"A8",
    X"09",X"00",X"04",X"08",X"04",X"00",X"21",X"21",
    X"00",X"FC",X"21",X"08",X"B7",X"00",X"C0",X"62",
    X"AA",X"00",X"04",X"00",X"B7",X"08",X"C0",X"7B",
    X"AA",X"04",X"FF",X"F7",X"00",X"C0",X"78",X"AA",
    X"00",X"FF",X"E7",X"00",X"C0",X"65",X"AA",X"04",
    X"00",X"04",X"08",X"04",X"01",X"00",X"00",X"00",
    X"FF",X"00",X"2A",X"FD",X"01",X"00",X"02",X"25",
    X"08",X"00",X"00",X"00",X"08",X"01",X"20",X"02",
    X"FD",X"00",X"00",X"F7",X"00",X"08",X"00",X"00",
    X"C0",X"28",X"FF",X"20",X"20",X"06",X"0F",X"21",
    X"00",X"20",X"02",X"FD",X"00",X"00",X"F6",X"FC",
    X"08",X"00",X"33",X"37",X"62",X"66",X"63",X"69",
    X"65",X"72",X"20",X"6F",X"61",X"78",X"75",X"58",
    X"20",X"20",X"20",X"20",X"20",X"00",X"20",X"69",
    X"69",X"72",X"00",X"20",X"64",X"6B",X"00",X"75",
    X"6E",X"68",X"69",X"20",X"20",X"64",X"66",X"41",
    X"61",X"64",X"73",X"78",X"54",X"69",X"63",X"20",
    X"63",X"6F",X"72",X"53",X"2E",X"20",X"79",X"73",
    X"74",X"2C",X"20",X"6B",X"0D",X"0A",X"64",X"20",
    X"74",X"0A",X"75",X"6F",X"69",X"20",X"20",X"64",
    X"66",X"41",X"66",X"20",X"74",X"69",X"69",X"0A",
    X"20",X"6E",X"66",X"6D",X"0A",X"73",X"67",X"65",
    X"69",X"66",X"20",X"69",X"74",X"63",X"6D",X"20",
    X"41",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );

-- This is a 16-bit SRAM split in 2 byte slices; so each slice will have two
-- bytes for each word of SRAM_SIZE
type t_sram is array(0 to SRAM_SIZE*2-1) of std_logic_vector(7 downto 0);
signal sram1 : t_sram := (
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );
signal sram0 : t_sram := (
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
    X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
    );

signal sram_chip_addr :     std_logic_vector(SRAM_ADDR_SIZE downto 1);
signal sram_output :        std_logic_vector(15 downto 0);

-- PROM table and interface signals --------------------------------------------

-- We'll simulate a 16-bit-wide static PROM (e.g. a Flash) with some serious
-- cycle time (70 or 90 ns).

constant PROM_SIZE : integer := 1024;
constant PROM_ADDR_SIZE : integer := log2(PROM_SIZE);

subtype t_prom_address is std_logic_vector(PROM_ADDR_SIZE-1 downto 0);
type t_prom is array(0 to PROM_SIZE-1) of t_word;

signal prom_rd_addr :       t_prom_address; 
signal prom_output :        std_logic_vector(7 downto 0);
signal prom_oe_n :          std_logic;

-- bram0 is LSB, bram3 is MSB
signal prom : t_prom := (
    X"3C04B000",X"24840154",X"0C000031",X"00000000",
    X"3C04B000",X"2484017D",X"0C000031",X"00000000",
    X"24080000",X"24090100",X"3C0A1234",X"354A5678",
    X"AD0A0000",X"21080004",X"214A0333",X"1D20FFFC",
    X"2129FFFF",X"24080000",X"24090100",X"3C0A1234",
    X"354A5678",X"3C0B1234",X"356B5678",X"8D0B0000",
    X"154B000A",X"21080004",X"214A0333",X"1D20FFFB",
    X"2129FFFF",X"3C04B000",X"248401BA",X"0C000031",
    X"00000000",X"08000027",X"00000000",X"3C04B000",
    X"248401BD",X"0C000031",X"00000000",X"3C04B000",
    X"248401C2",X"0C000031",X"00000000",X"3C04B000",
    X"2484019B",X"0C000031",X"00000000",X"0800002F",
    X"00000000",X"3C062000",X"80820000",X"10400008",
    X"24840001",X"8CC30020",X"30630002",X"1060FFFD",
    X"00000000",X"ACC20000",X"1000FFF7",X"00000000",
    X"03E00008",X"00000000",X"3C062000",X"3C07B000",
    X"24E70144",X"20A5FFFF",X"00A52820",X"00A52820",
    X"00A41006",X"3042000F",X"00E29021",X"82420000",
    X"8CC30020",X"30630002",X"1060FFFD",X"00000000",
    X"ACC20000",X"14A0FFF6",X"20A5FFFC",X"03E00008",
    X"00000000",X"30313233",X"34353637",X"38396162",
    X"63646566",X"0A0D4E6F",X"77207275",X"6E6E696E",
    X"67206672",X"6F6D2038",X"2D626974",X"20737461",
    X"74696320",X"6D656D6F",X"72790A0D",X"00546573",
    X"74696E67",X"2031362D",X"62697420",X"73746174",
    X"69632052",X"2F572E2E",X"2E200045",X"6E64206F",
    X"66207465",X"73742C20",X"70726F67",X"72616D20",
    X"66726F7A",X"656E2E0A",X"0D004F4B",X"00464149",
    X"4C000A0D",X"00202000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000"
    );



-- I/O devices -----------------------------------------------------------------

signal data_uart :          std_logic_vector(31 downto 0);
signal data_uart_status :   std_logic_vector(31 downto 0);
signal uart_tx_rdy :        std_logic := '1';
signal uart_rx_rdy :        std_logic := '1';

--------------------------------------------------------------------------------

signal clk :                std_logic := '0';
signal reset :              std_logic := '1';
signal interrupt :          std_logic := '0';
signal done :               std_logic := '0';

-- interface to asynchronous 16-bit-wide external SRAM
signal sram_address :       std_logic_vector(31 downto 0);
signal sram_data_rd :       std_logic_vector(15 downto 0);
signal sram_data_wr :       std_logic_vector(15 downto 0);
signal sram_byte_we_n :     std_logic_vector(1 downto 0);
signal sram_oe_n :          std_logic;

-- interface cpu-cache
signal cpu_data_addr :      t_word;
signal cpu_data_rd_vma :    std_logic;
signal cpu_data_rd :        t_word;
signal cpu_code_rd_addr :   t_pc;
signal cpu_code_rd :        t_word;
signal cpu_code_rd_vma :    std_logic;
signal cpu_data_wr :        t_word;
signal cpu_byte_we :        std_logic_vector(3 downto 0);
signal cpu_mem_wait :       std_logic;
signal cpu_ic_invalidate :  std_logic;
signal cpu_cache_enable :   std_logic;

-- interface to i/o
signal io_rd_data :         std_logic_vector(31 downto 0);
signal io_wr_data :         std_logic_vector(31 downto 0);
signal io_rd_addr :         std_logic_vector(31 downto 2);
signal io_wr_addr :         std_logic_vector(31 downto 2);
signal io_rd_vma :          std_logic;
signal io_byte_we :         std_logic_vector(3 downto 0);


--------------------------------------------------------------------------------
-- Logging signals


-- Log file
file log_file: TEXT open write_mode is "hw_sim_log.txt";

-- Console output log file
file con_file: TEXT open write_mode is "hw_sim_console_log.txt";

-- Maximum line size of for console output log. Lines longer than this will be
-- truncated.
constant CONSOLE_LOG_LINE_SIZE : integer := 1024*4;

-- Console log line buffer
signal con_line_buf :       string(1 to CONSOLE_LOG_LINE_SIZE);
signal con_line_ix :        integer := 1;

signal log_info :           t_log_info;

-- Debug signals ---------------------------------------------------------------


signal full_rd_addr :       std_logic_vector(31 downto 0);
signal full_wr_addr :       std_logic_vector(31 downto 0);
signal full_code_addr :     std_logic_vector(31 downto 0);


begin

    cpu: entity work.mips_cpu
    port map (
        interrupt   => '0',
        
        data_addr   => cpu_data_addr,
        data_rd_vma => cpu_data_rd_vma,
        data_rd     => cpu_data_rd,
        
        code_rd_addr=> cpu_code_rd_addr,
        code_rd     => cpu_code_rd,
        code_rd_vma => cpu_code_rd_vma,
        
        data_wr     => cpu_data_wr,
        byte_we     => cpu_byte_we,

        mem_wait    => cpu_mem_wait,
        cache_enable=> cpu_cache_enable,
        ic_invalidate=>cpu_ic_invalidate,
        
        clk         => clk,
        reset       => reset
    );


    cache: entity work.mips_cache
    generic map (
        BRAM_ADDR_SIZE => BRAM_ADDR_SIZE,
        SRAM_ADDR_SIZE => 32,-- we need the full address to decode sram vs flash
        LINE_SIZE =>      4,
        CACHE_SIZE =>     256
    )
    port map (
        clk             => clk,
        reset           => reset,
        
        -- Interface to CPU core
        data_addr       => cpu_data_addr,
        data_rd         => cpu_data_rd,
        data_rd_vma     => cpu_data_rd_vma,
                        
        code_rd_addr    => cpu_code_rd_addr,
        code_rd         => cpu_code_rd,
        code_rd_vma     => cpu_code_rd_vma,

        byte_we         => cpu_byte_we,
        data_wr         => cpu_data_wr,
                        
        mem_wait        => cpu_mem_wait,
        cache_enable    => cpu_cache_enable,
        ic_invalidate   => cpu_ic_invalidate,
        
        -- interface to FPGA i/o devices
        io_rd_data      => io_rd_data,
        io_wr_data      => io_wr_data,
        io_rd_addr      => io_rd_addr,
        io_wr_addr      => io_wr_addr,
        io_rd_vma       => io_rd_vma,
        io_byte_we      => io_byte_we,

        -- interface to synchronous 32-bit-wide FPGA BRAM
        bram_rd_data    => bram_rd_data,
        bram_wr_data    => bram_wr_data,
        bram_rd_addr    => bram_rd_addr,
        bram_wr_addr    => bram_wr_addr,
        bram_byte_we    => bram_byte_we,
        bram_data_rd_vma=> bram_data_rd_vma,
        
        -- interface to asynchronous 16-bit-wide external SRAM
        sram_address    => sram_address,
        sram_data_rd    => sram_data_rd,
        sram_data_wr    => sram_data_wr,
        sram_byte_we_n  => sram_byte_we_n,
        sram_oe_n       => sram_oe_n
    );

    ---------------------------------------------------------------------------
    -- Master clock: free running clock used as main module clock
    run_master_clock:
    process(done, clk)
    begin
        if done = '0' then
            clk <= not clk after T/2;
        end if;
    end process run_master_clock;

    drive_uut:
    process
    variable l : line;
    begin
        wait for T*4;
        reset <= '0';
        
        wait for T*SIMULATION_LENGTH;

        -- Flush console output to log console file (in case the end of the
        -- simulation caugh an unterminated line in the buffer)
        if con_line_ix > 1 then
            write(l, con_line_buf(1 to con_line_ix));
            writeline(con_file, l);
        end if;

        print("TB0 finished");
        done <= '1';
        wait;
        
    end process drive_uut;

    full_rd_addr <= cpu_data_addr;
    full_wr_addr <= cpu_data_addr(31 downto 2) & "00";
    full_code_addr <= cpu_code_rd_addr & "00";

    data_ram_block:
    process(clk)
    begin
        if clk'event and clk='1' then
            if reset='0' then
                bram_rd_data <= 
                    bram3(conv_integer(unsigned(bram_rd_addr))) &
                    bram2(conv_integer(unsigned(bram_rd_addr))) &
                    bram1(conv_integer(unsigned(bram_rd_addr))) &
                    bram0(conv_integer(unsigned(bram_rd_addr)));
                
                if bram_byte_we(3)='1' then
                    bram3(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr(31 downto 24);
                end if;
                if bram_byte_we(2)='1' then
                    bram2(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr(23 downto 16);
                end if;
                if bram_byte_we(1)='1' then
                    bram1(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr(15 downto  8);
                end if;
                if bram_byte_we(0)='1' then
                    bram0(conv_integer(unsigned(bram_wr_addr))) <= cpu_data_wr( 7 downto  0);
                end if;
            end if;
        end if;
    end process data_ram_block;

    sram_data_rd <= 
        X"00" & prom_output when sram_address(31 downto 27)="10110" else
        sram_output;
            


    -- Do a very basic simulation of an external SRAM ---------------

    sram_chip_addr <= sram_address(SRAM_ADDR_SIZE downto 1);

    -- FIXME should add some verification of /WE 
    sram_output <=
        sram1(conv_integer(unsigned(sram_chip_addr))) &
        sram0(conv_integer(unsigned(sram_chip_addr)))   when sram_oe_n='0'
        else (others => 'Z');

    simulated_sram_write:
    process(sram_byte_we_n, sram_address, sram_oe_n)
    begin
        -- Write cycle
        -- FIXME should add OE\ to write control logic
        if sram_byte_we_n'event or sram_address'event then
            if sram_byte_we_n(1)='0' then
                sram1(conv_integer(unsigned(sram_chip_addr))) <= sram_data_wr(15 downto  8);
            end if;
            if sram_byte_we_n(0)='0' then
                sram0(conv_integer(unsigned(sram_chip_addr))) <= sram_data_wr( 7 downto  0);
            end if;            
        end if;
    end process simulated_sram_write;


    -- Do a very basic simulation of an external PROM wired to the same bus 
    -- as the sram (both are static).
    
    prom_rd_addr <= sram_address(PROM_ADDR_SIZE+1 downto 2);
    
    prom_oe_n <= sram_oe_n;
    
    prom_output <=
        prom(conv_integer(unsigned(prom_rd_addr)))(31 downto 24) when prom_oe_n='0' and sram_address(1 downto 0)="00" else
        prom(conv_integer(unsigned(prom_rd_addr)))(23 downto 16) when prom_oe_n='0' and sram_address(1 downto 0)="01" else
        prom(conv_integer(unsigned(prom_rd_addr)))(15 downto  8) when prom_oe_n='0' and sram_address(1 downto 0)="10" else
        prom(conv_integer(unsigned(prom_rd_addr)))( 7 downto  0) when prom_oe_n='0' and sram_address(1 downto 0)="11" else
        (others => 'Z');
    
    
    simulated_io:
    process(clk)
    variable i : integer;
    variable uart_data : integer;
    begin
        if clk'event and clk='1' then
            
            if io_byte_we/="0000" then
                if io_wr_addr(31 downto 28)=X"2" then
                    -- Write to UART
                    
                    -- If we're simulating the UART TX time, pulse RDY low
                    if SIMULATED_UART_TX_TIME > 0 us then
                        uart_tx_rdy <= '0', '1' after SIMULATED_UART_TX_TIME;
                    end if;
                    
                    -- TX data may come from the high or low byte (opcodes.s
                    -- uses high byte, no_op.c uses low)
                    if io_byte_we(0)='1' then
                        uart_data := conv_integer(unsigned(io_wr_data(7 downto 0)));
                    else
                        uart_data := conv_integer(unsigned(io_wr_data(31 downto 24)));
                    end if;
                    
                    -- UART TX data goes to output after a bit of line-buffering
                    -- and editing
                    if uart_data = 10 then
                        -- CR received: print output string and clear it
                        print(con_file, con_line_buf(1 to con_line_ix));
                        con_line_ix <= 1;
                        for i in 1 to con_line_buf'high loop
                           con_line_buf(i) <= ' ';
                        end loop;
                    elsif uart_data = 13 then
                        -- ignore LF
                    else
                        -- append char to output string
                        if con_line_ix < con_line_buf'high then
                            con_line_buf(con_line_ix) <= character'val(uart_data);
                            con_line_ix <= con_line_ix + 1;
                        end if;
                    end if;
                end if;
            end if;
        end if;
    end process simulated_io;

    -- UART read registers; only status, and hardwired, for the time being
    io_rd_data <= X"00000003";
    data_uart <= data_uart_status;
    data_uart_status <= X"0000000" & "00" & uart_tx_rdy & uart_rx_rdy;

    log_execution:
    process
    begin
        log_cpu_activity(clk, reset, done, 
                         "mips_tb2/cpu", log_info, "log_info", 
                         X"BFC00000", log_file);
        wait;
    end process log_execution;

    
end architecture testbench;
