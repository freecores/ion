--------------------------------------------------------------------------------
-- File built automatically for project 'Hello World' by bin2hdl.py
--------------------------------------------------------------------------------
-- Synthesizable ROM implemented on regular FPGA BLock RAM MPU.
--
-- Meant to be used as bootstrap code ROM in project ION, hence the fixed
-- entity name.
--
-- This package provides constants and types that will be used wherever the code
-- BRAM is implemented, presumably in the mips_mpu module (see that module for
-- an usage example).
--
-- Note that no vendor-specific stuff needs to be used at all to infer the
-- read-only, single port BRAM we're interested in.
--------------------------------------------------------------------------------
-- Copyright (C) 2011 Jose A. Ruiz
--                                                              
-- This source file may be used and distributed without         
-- restriction provided that this copyright statement is not    
-- removed from the file and that any derivative work contains  
-- the original copyright notice and the associated disclaimer. 
--                                                              
-- This source file is free software; you can redistribute it   
-- and/or modify it under the terms of the GNU Lesser General   
-- Public License as published by the Free Software Foundation; 
-- either version 2.1 of the License, or (at your option) any   
-- later version.                                               
--                                                              
-- This source is distributed in the hope that it will be       
-- useful, but WITHOUT ANY WARRANTY; without even the implied   
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      
-- PURPOSE.  See the GNU Lesser General Public License for more 
-- details.                                                     
--                                                              
-- You should have received a copy of the GNU Lesser General    
-- Public License along with this source; if not, download it   
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mips_pkg.all;

package code_rom_pkg is

-- BRAM table and address word sizes...
constant CODE_BRAM_SIZE : integer := 2048;
constant CODE_BRAM_ADDR_SIZE : integer := log2(CODE_BRAM_SIZE);
subtype t_bram_address is std_logic_vector(CODE_BRAM_ADDR_SIZE-1 downto 0);
-- ...and the type of the actual table that will hold the data.
type t_bram is array(0 to (CODE_BRAM_SIZE)-1) of t_word;

-- This constant defines the contents of the BRAM.
constant code_bram :                  t_bram := (
    X"1000007C",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"401A6800",X"001AD082",X"335A001F",X"341B0008",
    X"135B0009",X"237B0001",X"135B0005",X"237B0001",
    X"175B0007",X"00000000",X"0BF000A2",X"00000000",
    X"0BF00072",X"00000000",X"0BF00072",X"00000000",
    X"0BF00072",X"00000000",X"401B7000",X"401A6800",
    X"001AD7C2",X"335A0001",X"17400003",X"237B0004",
    X"03600008",X"00000000",X"237B0004",X"03600008",
    X"42000010",X"40046000",X"3084FFFE",X"40846000",
    X"0FF00086",X"00000000",X"3C04BFC0",X"248406B4",
    X"00800008",X"00000000",X"3C050001",X"40046000",
    X"3084FFFF",X"00852825",X"40856000",X"24040000",
    X"24060000",X"240500FF",X"AC860000",X"00C5082A",
    X"1420FFFD",X"20C60001",X"24040000",X"24060000",
    X"240500FF",X"8C800000",X"20840010",X"00C5082A",
    X"1420FFFC",X"20C60001",X"3C050002",X"40046000",
    X"3084FFFF",X"00852825",X"03E00008",X"40856000",
    X"00000000",X"00000000",X"3C1B0000",X"277B003C",
    X"AF7DFFF0",X"AF7FFFEC",X"AF68FFE8",X"AF69FFE4",
    X"AF6AFFE0",X"0360E821",X"40087000",X"8D1A0000",
    X"401B6800",X"0770002D",X"00000000",X"001A4E82",
    X"3928001F",X"1100001F",X"3928001C",X"11000013",
    X"00000000",X"3C082001",X"AD1A0400",X"8FAAFFE0",
    X"8FA9FFE4",X"8FA8FFE8",X"8FBFFFEC",X"8FBDFFF0",
    X"401B7000",X"401A6800",X"001AD7C2",X"335A0001",
    X"17400003",X"237B0004",X"03600008",X"00000000",
    X"237B0004",X"03600008",X"42000010",X"335B003F",
    X"3B680020",X"11000014",X"3B680021",X"1100001C",
    X"00000000",X"3C082001",X"AD1A0400",X"0BF000B7",
    X"00000000",X"335B003F",X"3B680000",X"1100001E",
    X"3B680004",X"11000029",X"00000000",X"3C082001",
    X"AD1A0400",X"0BF000B7",X"00000000",X"8D1A0004",
    X"03E00008",X"00000000",X"0FF00161",X"3C0A8000",
    X"00004021",X"036A4824",X"15200003",X"000A5042",
    X"1540FFFC",X"25080001",X"0BF00117",X"0100D821",
    X"0FF00161",X"3C0A8000",X"00004021",X"036A4824",
    X"11200003",X"000A5042",X"1540FFFC",X"25080001",
    X"0BF00117",X"0100D821",X"0FF00161",X"00000000",
    X"001A4182",X"3108001F",X"001A4AC2",X"3129001F",
    X"01095021",X"000A5023",X"254A001F",X"015BD804",
    X"015BD806",X"0BF00117",X"011BD806",X"0FF00161",
    X"00000000",X"001A4182",X"3108001F",X"001A4AC2",
    X"3129001F",X"01284823",X"00095823",X"256B001F",
    X"011B4804",X"3C0AFFFF",X"354AFFFF",X"016A5004",
    X"016A5006",X"010A5004",X"012A4824",X"01405027",
    X"0FF00161",X"001AD140",X"001AD142",X"036AD824",
    X"0369D825",X"0BF00117",X"00000000",X"001A4C02",
    X"3129001F",X"3C08BFC0",X"25080484",X"000948C0",
    X"01094020",X"01000008",X"00000000",X"0BF000B7",
    X"00000000",X"0BF0011F",X"37600000",X"0BF0011F",
    X"37610000",X"0BF0011F",X"37620000",X"0BF0011F",
    X"37630000",X"0BF0011F",X"37640000",X"0BF0011F",
    X"37650000",X"0BF0011F",X"37660000",X"0BF0011F",
    X"37670000",X"0BF0011F",X"AFBBFFE8",X"0BF0011F",
    X"AFBBFFE4",X"0BF0011F",X"AFBBFFE0",X"0BF0011F",
    X"376B0000",X"0BF0011F",X"376C0000",X"0BF0011F",
    X"376D0000",X"0BF0011F",X"376E0000",X"0BF0011F",
    X"376F0000",X"0BF0011F",X"37700000",X"0BF0011F",
    X"37710000",X"0BF0011F",X"37720000",X"0BF0011F",
    X"37730000",X"0BF0011F",X"37740000",X"0BF0011F",
    X"37750000",X"0BF0011F",X"37760000",X"0BF0011F",
    X"37770000",X"0BF0011F",X"37780000",X"0BF0011F",
    X"37790000",X"0BF0011F",X"377A0000",X"0BF0011F",
    X"377B0000",X"0BF0011F",X"377C0000",X"0BF0011F",
    X"AFBBFFEC",X"0BF0011F",X"377E0000",X"0BF0011F",
    X"AFBBFFF0",X"AFBF0000",X"001ADD42",X"337B001F",
    X"3C08BFC0",X"250805B4",X"001BD8C0",X"011B4020",
    X"0100F809",X"00000000",X"8FBF0000",X"03E00008",
    X"00000000",X"03E00008",X"341B0000",X"03E00008",
    X"343B0000",X"03E00008",X"345B0000",X"03E00008",
    X"347B0000",X"03E00008",X"349B0000",X"03E00008",
    X"34BB0000",X"03E00008",X"34DB0000",X"03E00008",
    X"34FB0000",X"03E00008",X"8FBBFFE8",X"03E00008",
    X"8FBBFFE4",X"03E00008",X"8FBBFFE0",X"03E00008",
    X"357B0000",X"03E00008",X"359B0000",X"03E00008",
    X"35BB0000",X"03E00008",X"35DB0000",X"03E00008",
    X"35FB0000",X"03E00008",X"361B0000",X"03E00008",
    X"363B0000",X"03E00008",X"365B0000",X"03E00008",
    X"367B0000",X"03E00008",X"369B0000",X"03E00008",
    X"36BB0000",X"03E00008",X"36DB0000",X"03E00008",
    X"36FB0000",X"03E00008",X"371B0000",X"03E00008",
    X"373B0000",X"03E00008",X"375B0000",X"03E00008",
    X"377B0000",X"03E00008",X"379A0000",X"03E00008",
    X"8FBBFFF0",X"03E00008",X"37DB0000",X"03E00008",
    X"8FBBFFEC",X"3C1C0000",X"279C7FF0",X"3C050000",
    X"24A50000",X"3C040000",X"24840000",X"3C1D0000",
    X"27BD0428",X"ACA00000",X"00A4182A",X"1460FFFD",
    X"24A50004",X"3C040000",X"24840000",X"3C05BFC0",
    X"24A50E60",X"10A4000B",X"00000000",X"3C100000",
    X"26100000",X"12000007",X"00000000",X"8CA80000",
    X"24A50004",X"AC880000",X"24840004",X"1600FFFB",
    X"2610FFFC",X"0FF001CD",X"00000000",X"0BF001CB",
    X"00000000",X"3C04BFC0",X"27BDFFE8",X"AFBF0014",
    X"0FF00340",X"24840E04",X"3C04BFC0",X"0FF00340",
    X"24840E2C",X"3C04BFC0",X"8FBF0014",X"24840E44",
    X"0BF00340",X"27BD0018",X"10800009",X"00000000",
    X"8C820000",X"00000000",X"A0450000",X"8C820000",
    X"00000000",X"24420001",X"03E00008",X"AC820000",
    X"0BF0036E",X"00A02021",X"27BDFFD8",X"AFB20018",
    X"AFB10014",X"AFB00010",X"AFBF0024",X"AFB40020",
    X"AFB3001C",X"00C09021",X"00808821",X"18C00032",
    X"00A08021",X"90A20000",X"00000000",X"1040003D",
    X"00A01021",X"00001821",X"24420001",X"90440000",
    X"00000000",X"1480FFFC",X"24630001",X"0072102A",
    X"14400002",X"02439023",X"00009021",X"30E20002",
    X"10400022",X"30E70001",X"10E00022",X"24140030",
    X"00009821",X"92050000",X"00000000",X"10A00008",
    X"00000000",X"02202021",X"0FF001DA",X"26100001",
    X"92050000",X"00000000",X"14A0FFFA",X"26730001",
    X"1A400008",X"02408021",X"2610FFFF",X"02202021",
    X"0FF001DA",X"02802821",X"1600FFFC",X"2610FFFF",
    X"02729821",X"8FBF0024",X"02601021",X"8FB40020",
    X"8FB3001C",X"8FB20018",X"8FB10014",X"8FB00010",
    X"03E00008",X"27BD0028",X"30E70001",X"14E0FFE0",
    X"24140020",X"1A40FFDE",X"02409821",X"2673FFFF",
    X"02202021",X"0FF001DA",X"02802821",X"1660FFFC",
    X"2673FFFF",X"26730001",X"02409821",X"0BF00205",
    X"00009021",X"00001821",X"0BF001FF",X"02439023",
    X"27BDFFC8",X"AFB40030",X"AFB20028",X"AFB10024",
    X"AFBF0034",X"AFB3002C",X"AFB00020",X"00A01021",
    X"8FB40048",X"8FB2004C",X"10A0003F",X"00808821",
    X"14E00031",X"2403000A",X"00003821",X"10400049",
    X"A3A0001B",X"8FA50050",X"27B3001B",X"24A5FFC6",
    X"14C00002",X"0046001B",X"0007000D",X"00001810",
    X"2864000A",X"00000000",X"14C00002",X"0046001B",
    X"0007000D",X"00001012",X"14800002",X"2673FFFF",
    X"00651821",X"24630030",X"1440FFF1",X"A2630000",
    X"14E00010",X"00000000",X"00008021",X"02202021",
    X"02602821",X"02803021",X"0FF001E6",X"02403821",
    X"8FBF0034",X"00501021",X"8FB40030",X"8FB3002C",
    X"8FB20028",X"8FB10024",X"8FB00020",X"03E00008",
    X"27BD0038",X"1280000F",X"32420002",X"1040000D",
    X"02202021",X"0FF001DA",X"2405002D",X"2694FFFF",
    X"0BF0025B",X"24100001",X"14C3FFD0",X"00003821",
    X"04A1FFCE",X"00000000",X"00051023",X"0BF00243",
    X"24070001",X"2673FFFF",X"2402002D",X"A2620000",
    X"0BF0025B",X"00008021",X"27A50010",X"02803021",
    X"02403821",X"24020030",X"A3A20010",X"0FF001E6",
    X"A3A00011",X"8FBF0034",X"8FB40030",X"8FB3002C",
    X"8FB20028",X"8FB10024",X"8FB00020",X"03E00008",
    X"27BD0038",X"10E0FFCC",X"27B3001B",X"0BF00269",
    X"00000000",X"27BDFFB8",X"AFB40038",X"AFB00028",
    X"AFBF0044",X"AFB60040",X"AFB5003C",X"AFB30034",
    X"AFB20030",X"AFB1002C",X"00A08021",X"90A50000",
    X"0080A021",X"10A000A0",X"AFA60050",X"00009021",
    X"24130025",X"2415002D",X"24110030",X"3C16BFC0",
    X"14B30053",X"00000000",X"26100001",X"92050000",
    X"00000000",X"10A0003E",X"00000000",X"10B3004C",
    X"00000000",X"10B50054",X"00000000",X"00001821",
    X"14B10007",X"24A2FFD0",X"26100001",X"92050000",
    X"00000000",X"10B1FFFC",X"34630002",X"24A2FFD0",
    X"304200FF",X"2C42000A",X"1040000D",X"00001021",
    X"00022040",X"000210C0",X"00821021",X"26100001",
    X"00451021",X"92050000",X"00000000",X"24A4FFD0",
    X"308400FF",X"2C84000A",X"1480FFF5",X"2442FFD0",
    X"24040073",X"10A4003C",X"24040064",X"10A40046",
    X"02802021",X"24040078",X"10A40051",X"02802021",
    X"24040058",X"10A40055",X"02802021",X"24040075",
    X"10A40060",X"02802021",X"24040063",X"14A40024",
    X"26100001",X"8FA90050",X"27A50020",X"8D280000",
    X"02802021",X"25290004",X"00403021",X"00603821",
    X"AFA90050",X"A3A80020",X"0FF001E6",X"A3A00021",
    X"92050000",X"00000000",X"14A0FFBD",X"02429021",
    X"12800004",X"00000000",X"8E820000",X"00000000",
    X"A0400000",X"8FBF0044",X"02401021",X"8FB60040",
    X"8FB5003C",X"8FB40038",X"8FB30034",X"8FB20030",
    X"8FB1002C",X"8FB00028",X"03E00008",X"27BD0048",
    X"0FF001DA",X"02802021",X"26520001",X"26100001",
    X"92050000",X"00000000",X"14A0FFA5",X"00000000",
    X"0BF002E8",X"00000000",X"26100001",X"92050000",
    X"0BF002B0",X"24030001",X"8FA40050",X"00000000",
    X"8C850000",X"24840004",X"10A00031",X"AFA40050",
    X"02802021",X"00403021",X"0FF001E6",X"00603821",
    X"0BF002FB",X"02429021",X"8FA80050",X"00000000",
    X"8D050000",X"2406000A",X"25080004",X"24070001",
    X"AFA20010",X"24020061",X"AFA80050",X"AFA30014",
    X"0FF00234",X"AFA20018",X"0BF002FB",X"02429021",
    X"8FA80050",X"00000000",X"8D050000",X"24060010",
    X"25080004",X"0BF00318",X"00003821",X"8FA80050",
    X"00000000",X"8D050000",X"24060010",X"25080004",
    X"AFA20010",X"00003821",X"24020041",X"AFA80050",
    X"AFA30014",X"0FF00234",X"AFA20018",X"0BF002FB",
    X"02429021",X"8FA80050",X"00000000",X"8D050000",
    X"2406000A",X"25080004",X"0BF00318",X"00003821",
    X"0BF0030C",X"26C50E58",X"0BF002E8",X"00009021",
    X"27BDFFE0",X"27A20024",X"00801821",X"AFA50024",
    X"AFA60028",X"00002021",X"00602821",X"00403021",
    X"AFBF001C",X"AFA7002C",X"0FF00291",X"AFA20010",
    X"8FBF001C",X"00000000",X"03E00008",X"27BD0020",
    X"27BDFFE0",X"27A20028",X"AFA40020",X"AFA60028",
    X"27A40020",X"00403021",X"AFBF001C",X"AFA7002C",
    X"0FF00291",X"AFA20010",X"8FBF001C",X"00000000",
    X"03E00008",X"27BD0020",X"27BDFFE0",X"27A2002C",
    X"AFA40020",X"00C02821",X"27A40020",X"00403021",
    X"AFBF001C",X"AFA7002C",X"0FF00291",X"AFA20010",
    X"8FBF001C",X"00000000",X"03E00008",X"27BD0020",
    X"03E00008",X"00001021",X"00801021",X"3C052000",
    X"8CA30020",X"00000000",X"30630002",X"1060FFFC",
    X"3C032000",X"AC620000",X"03E00008",X"00000000",
    X"3C032000",X"8C620020",X"00000000",X"30420001",
    X"1040FFFC",X"3C022000",X"8C420000",X"03E00008",
    X"00021602",X"636F6D70",X"696C6520",X"74696D65",
    X"3A204A75",X"6E202038",X"20323031",X"32202D2D",
    X"2032333A",X"30343A32",X"360A0000",X"67636320",
    X"76657273",X"696F6E3A",X"2020342E",X"352E320A",
    X"00000000",X"0A0A4865",X"6C6C6F20",X"576F726C",
    X"64210A0A",X"0A000000",X"286E756C",X"6C290000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000",
    X"00000000",X"00000000",X"00000000",X"00000000"
    );

end package;
